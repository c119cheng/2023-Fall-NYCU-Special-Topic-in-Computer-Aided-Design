module c10000 (I4737, I4052, I3510, I389, I2768, I29, I1544, I1759, I1646, I4182, I4743, I4001, I2233, I397, I425, I1494, I2103, I2521, I1222, I491, I1594, I900, I4728, I3598, I1718, I3047, I2709, I4555, I4806, I2484, I193, I4557, I3044, I2462, I192, I2748, I4692, I1021, I16, I282, I1699, I3402, I3118, I2732, I3270, I2113, I76, I2613, I1430, I3071, I1076, I2564, I915, I1601, I391, I2780, I379, I1870, I334, I1769, I4135, I2866, I4047, I4323, I1347, I3300, I1930, I3395, I2693, I3699, I2725, I3560, I4190, I4657, I1631, I3694, I2002, I815, I4439, I3306, I1977, I4928, I523, I2073, I4846, I3473, I4290, I3949, I4983, I736, I4109, I604, I559, I2735, I3152, I3700, I3372, I832, I3570, I767, I4835, I2086, I1840, I2785, I2666, I3575, I721, I4665, I417, I69, I3588, I1052, I2624, I422, I875, I817, I500, I3534, I766, I67, I534, I1185, I4594, I3781, I3009, I2094, I1410, I989, I1257, I2065, I4359, I3100, I22, I3973, I1237, I328, I1662, I848, I3684, I1447, I2675, I1230, I2378, I392, I1738, I4152, I3989, I242, I778, I2389, I2022, I1561, I3968, I2097, I3098, I2004, I555, I1099, I2117, I4272, I1203, I2154, I4626, I4891, I4481, I4220, I600, I2811, I2343, I4568, I1876, I2418, I4035, I458, I1775, I3696, I3379, I4391, I3942, I1233, I4711, I925, I2059, I1563, I3892, I4287, I686, I4645, I12, I754, I3654, I526, I4102, I1665, I408, I1771, I2043, I1479, I677, I226, I154, I3540, I1551, I4076, I2514, I587, I4773, I800, I4575, I3688, I2492, I3773, I4549, I4824, I4795, I4628, I77, I568, I2125, I1816, I1355, I4260, I2376, I2581, I513, I2013, I339, I691, I2929, I1654, I271, I2582, I3440, I3791, I774, I3444, I1461, I1024, I2177, I4176, I3660, I1379, I4432, I1781, I346, I1323, I3459, I1117, I4934, I1317, I2480, I4904, I3151, I2409, I3380, I2758, I2118, I4145, I3464, I1256, I197, I3414, I2734, I808, I775, I1285, I2280, I1420, I1463, I3134, I1393, I1900, I4156, I3256, I1426, I739, I3442, I997, I2927, I1831, I3852, I4357, I57, I2353, I3358, I4171, I906, I3627, I1627, I119, I2036, I1815, I4049, I1482, I1079, I2744, I3809, I63, I635, I3648, I2070, I1574, I1155, I3638, I3235, I4378, I4048, I764, I4101, I3333, I1440, I4590, I2267, I3906, I4057, I3879, I2106, I2179, I914, I3900, I2241, I4334, I2061, I3512, I2447, I2095, I1637, I3361, I369, I521, I2683, I1097, I1301, I3172, I1597, I1659, I4160, I2777, I3480, I859, I58, I4023, I913, I3777, I3317, I2202, I2659, I3636, I4079, I493, I4195, I443, I678, I3110, I3750, I208, I599, I3966, I2437, I1992, I2152, I2828, I1877, I1540, I4883, I2033, I1160, I3324, I4763, I2702, I1617, I3673, I2713, I4255, I239, I1572, I2146, I1826, I4546, I4243, I948, I306, I3943, I3025, I1473, I1335, I2458, I4392, I2743, I3720, I4879, I821, I2865, I1522, I4856, I991, I2433, I3817, I1418, I2032, I1863, I74, I1966, I4944, I1116, I4054, I2160, I3722, I620, I418, I2137, I4394, I1140, I3345, I2475, I2224, I1896, I1260, I3215, I3065, I3058, I2988, I1553, I3077, I2364, I2769, I2450, I1204, I3138, I1868, I2868, I4573, I1320, I3237, I3656, I3602, I3326, I2588, I4234, I4369, I4646, I3406, I2642, I950, I3936, I1353, I1867, I1899, I4332, I4119, I2121, I3893, I3188, I1382, I1383, I3719, I623, I3170, I2162, I3164, I742, I1327, I2861, I1223, I1298, I4129, I2906, I2093, I4146, I4343, I1488, I1096, I4844, I969, I1330, I4830, I1710, I3316, I4804, I3026, I2392, I4469, I176, I918, I2858, I4405, I148, I3198, I240, I497, I2691, I856, I331, I1409, I3577, I3523, I2503, I510, I3457, I4760, I1112, I4571, I1108, I1915, I977, I585, I3780, I3296, I3815, I18, I5, I3297, I1190, I2937, I3663, I1265, I3017, I1004, I3771, I2217, I3054, I4285, I1492, I4649, I2049, I1073, I4601, I2633, I3685, I3181, I4624, I3935, I929, I2647, I4110, I2730, I905, I3806, I4616, I1683, I2368, I4225, I332, I1679, I720, I2677, I95, I90, I1857, I1487, I227, I1752, I19, I1425, I400, I575, I3192, I2188, I3066, I2427, I2425, I3216, I2003, I695, I1817, I4120, I2112, I1, I4261, I3969, I71, I553, I3996, I3325, I4370, I586, I3328, I3513, I1811, I4655, I1307, I3488, I1229, I3231, I3413, I1061, I3617, I3162, I3336, I2222, I4630, I3782, I499, I4203, I1321, I1660, I312, I3521, I2416, I2303, I1792, I2635, I3346, I155, I3376, I842, I4933, I3839, I3576, I3353, I698, I4526, I970, I3059, I4041, I4075, I2213, I2272, I2903, I4714, I4751, I4371, I3661, I3301, I433, I96, I2957, I3863, I477, I1159, I713, I1325, I1034, I1842, I2540, I3185, I4324, I4467, I70, I380, I610, I1132, I1694, I2193, I1465, I4602, I2109, I2099, I179, I243, I4447, I1178, I3946, I3896, I2216, I2127, I1514, I954, I1127, I3284, I4200, I4674, I3020, I4515, I4828, I2438, I3561, I214, I782, I1963, I2697, I3165, I4910, I2576, I2051, I858, I1768, I2688, I1936, I2225, I2523, I4545, I2789, I3396, I703, I1750, I2435, I471, I1029, I876, I4956, I3496, I2373, I1645, I4294, I1311, I267, I786, I2479, I2145, I228, I4621, I451, I1496, I1834, I4690, I206, I3472, I464, I4745, I2722, I980, I934, I2834, I3486, I1081, I1794, I1349, I4873, I2573, I2682, I4163, I78, I4331, I4045, I1384, I631, I868, I4902, I4963, I1648, I1879, I2044, I3934, I3708, I3425, I3903, I1415, I2305, I606, I2965, I2947, I196, I4169, I4942, I3200, I4524, I3793, I3668, I1669, I2676, I4158, I4787, I3349, I3417, I2251, I4863, I2180, I4142, I440, I1240, I3535, I2342, I2481, I59, I1143, I1974, I2219, I1859, I191, I897, I1247, I1451, I4778, I4868, I3386, I2223, I2601, I3869, I1677, I3153, I4679, I845, I829, I1017, I4382, I662, I1853, I676, I1972, I820, I3659, I3904, I1546, I4148, I447, I185, I313, I2765, I1839, I2348, I2312, I244, I2337, I4066, I1557, I3115, I3508, I2547, I2369, I603, I3147, I1692, I2815, I3778, I1345, I3236, I1386, I3178, I2358, I27, I2388, I3243, I1071, I382, I756, I87, I4821, I2108, I3429, I890, I4409, I1716, I3203, I4880, I1777, I4849, I1368, I1068, I1422, I3929, I3280, I349, I2083, I4799, I3323, I4980, I588, I2706, I3649, I4161, I2028, I4666, I365, I1477, I3040, I709, I4107, I1395, I479, I1552, I1957, I1709, I355, I803, I4730, I1605, I120, I990, I573, I2962, I921, I4346, I3878, I1953, I2453, I2580, I386, I4712, I2354, I2570, I4112, I4976, I4802, I4611, I2849, I1157, I3538, I3850, I3703, I51, I3202, I4710, I2895, I2796, I4012, I1293, I4221, I1003, I3201, I1455, I784, I4689, I2907, I4259, I2993, I1333, I4192, I2627, I4936, I2471, I177, I2830, I3584, I2585, I2641, I3171, I1567, I1517, I2631, I580, I115, I1770, I2363, I1556, I3279, I2140, I2669, I3272, I3639, I292, I3907, I735, I4991, I2824, I4913, I3594, I3503, I1991, I1761, I2994, I3796, I509, I241, I3415, I3435, I2211, I4958, I1723, I1043, I931, I4619, I152, I3299, I3046, I2417, I1790, I3759, I3601, I4410, I2075, I34, I54, I325, I4924, I1401, I1721, I2320, I1458, I939, I219, I2339, I750, I3334, I2421, I3108, I1988, I1469, I2276, I2428, I1365, I3772, I3365, I1454, I2512, I4486, I3391, I1039, I4808, I2201, I2087, I3183, I4859, I1032, I565, I4170, I4473, I2716, I3739, I4452, I3976, I1596, I2472, I1524, I3860, I4113, I3458, I1907, I1255, I3669, I3580, I3536, I1805, I4961, I622, I2609, I1188, I4300, I412, I1622, I3155, I1057, I7, I1405, I935, I2727, I2129, I1955, I968, I4459, I891, I641, I1516, I1388, I757, I715, I1727, I2749, I4062, I3479, I2525, I2754, I3314, I250, I4815, I4199, I8, I1786, I225, I4803, I3619, I124, I362, I2517, I2872, I569, I402, I3775, I618, I4845, I3304, I4987, I1528, I1909, I996, I855, I539, I1212, I494, I722, I4684, I4698, I4886, I1176, I4926, I3651, I4027, I912, I4599, I1197, I321, I2753, I4464, I1022, I4030, I1693, I1643, I3836, I4905, I780, I490, I2586, I1119, I4217, I4542, I3160, I2707, I3266, I2150, I4328, I4484, I3578, I2327, I1600, I3798, I3705, I984, I1196, I3094, I3339, I4927, I2394, I3123, I3606, I694, I3103, I1880, I3667, I822, I2237, I305, I903, I4201, I4028, I2157, I1030, I1241, I644, I4282, I3554, I4850, I1090, I1098, I1436, I1765, I1827, I4291, I2680, I3792, I295, I3456, I3455, I3840, I3449, I4676, I3611, I4785, I702, I4925, I2290, I118, I704, I1807, I3928, I1089, I1226, I1216, I4126, I828, I3029, I3811, I577, I3484, I272, I1838, I4986, I3310, I3672, I144, I2531, I4695, I4111, I3709, I3366, I3438, I2166, I1576, I1134, I4884, I3268, I3149, I661, I4015, I3991, I1999, I4615, I3374, I4185, I3820, I2460, I2257, I4985, I2701, I4607, I2473, I1446, I1141, I81, I2203, I4007, I3393, I4513, I2287, I2419, I3559, I1939, I2893, I1381, I4056, I275, I4860, I1829, I2920, I262, I1168, I4578, I4356, I4437, I2430, I3533, I1296, I3988, I765, I3671, I3910, I4984, I4982, I4092, I2714, I1798, I104, I3193, I4498, I431, I264, I291, I3079, I3564, I2837, I4000, I2040, I1731, I1923, I2597, I310, I4544, I3514, I2846, I3628, I1315, I399, I1045, I546, I3050, I411, I3221, I1932, I1352, I2165, I3282, I1856, I1075, I2314, I790, I4400, I372, I435, I1890, I2014, I1394, I1275, I1527, I1470, I2844, I4496, I4857, I2221, I3827, I4438, I2956, I3916, I2311, I3692, I4070, I3116, I4264, I2578, I4506, I3359, I1545, I974, I4805, I3757, I3468, I1067, I2739, I3209, I2829, I4068, I4069, I456, I3142, I602, I198, I4890, I290, I358, I4969, I4648, I2850, I1059, I2139, I3084, I3995, I2069, I3971, I1566, I1541, I3641, I1308, I1613, I578, I2919, I3812, I692, I3873, I1931, I315, I1326, I4222, I3360, I3315, I2562, I3001, I186, I461, I2301, I2340, I3506, I3052, I793, I4389, I4197, I2604, I288, I684, I3591, I2254, I663, I1933, I2658, I2720, I1390, I2784, I2657, I3061, I232, I48, I1306, I2831, I937, I1644, I2309, I4304, I888, I1614, I3545, I3717, I4297, I3765, I252, I4522, I13, I1148, I453, I2077, I1580, I4050, I478, I1642, I792, I1336, I2974, I4008, I3822, I3888, I3630, I3060, I4417, I4640, I728, I1700, I814, I4210, I1086, I1364, I238, I2493, I4764, I4653, I2068, I220, I3593, I2400, I3056, I567, I3992, I1400, I4771, I1942, I933, I2605, I4096, I1149, I1016, I4885, I2296, I1995, I2989, I1658, I2238, I3122, I1267, I1284, I1290, I4211, I3653, I690, I1742, I904, I1146, I1799, I4783, I2035, I2515, I3861, I343, I2482, I2380, I1785, I4431, I2352, I2005, I3608, I1575, I404, I3932, I165, I133, I256, I1421, I4011, I1123, I341, I1033, I4719, I3481, I960, I883, I2101, I1782, I2334, I3970, I1125, I2198, I167, I819, I2134, I4669, I2574, I3712, I518, I2971, I4822, I4471, I4660, I4322, I3062, I992, I1866, I1773, I3015, I2662, I3530, I2026, I1864, I3168, I854, I4420, I79, I1702, I2274, I2909, I3944, I4915, I64, I2606, I2857, I347, I4298, I1489, I3963, I4734, I3416, I4277, I2148, I2361, I345, I4336, I4033, I3662, I2478, I3981, I1434, I2596, I2779, I388, I2090, I4548, I2273, I3931, I4659, I2260, I572, I1506, I1485, I3180, I4177, I2483, I1371, I3163, I2817, I4078, I2835, I1847, I1937, I4407, I2924, I189, I4570, I1951, I4465, I1445, I3232, I711, I4629, I4931, I273, I4038, I871, I2381, I1595, I2391, I4143, I3629, I172, I92, I1439, I2345, I3565, I863, I732, I3568, I1173, I3408, I3832, I4532, I1103, I4319, I3621, I670, I314, I4869, I2042, I4091, I3214, I3248, I4090, I444, I432, I3704, I551, I2818, I3738, I25, I1889, I1500, I4635, I2900, I446, I336, I2102, I615, I4762, I3397, I983, I2175, I3625, I212, I956, I1640, I2133, I2184, I169, I4838, I4789, I2944, I2300, I3918, I3616, I1929, I1239, I1818, I4966, I2958, I2612, I1904, I3657, I1292, I4348, I2485, I1878, I2859, I741, I1536, I4114, I570, I1959, I3899, I4625, I761, I3724, I1970, I4269, I1869, I353, I4862, I257, I1862, I492, I2474, I4576, I1590, I795, I1823, I3961, I1664, I2788, I2724, I4306, I1350, I1641, I919, I4002, I4493, I1726, I2465, I650, I2250, I1996, I1219, I4579, I1402, I4800, I3876, I1391, I4016, I561, I2147, I1309, I3362, I1633, I1751, I3557, I3945, I743, I213, I1162, I455, I1753, I3953, I3491, I2856, I3341, I4807, I594, I3956, I3562, I2092, I3068, I503, I108, I2350, I4643, I2464, I1051, I2904, I41, I396, I483, I4031, I3392, I3294, I853, I4779, I2726, I23, I164, I2534, I139, I2397, I4131, I2404, I2046, I3154, I665, I4833, I957, I1011, I1908, I2072, I745, I520, I3891, I1107, I1289, I1533, I2420, I2731, I2151, I3027, I4067, I877, I697, I4748, I126, I4775, I3810, I1571, I3537, I4208, I3319, I3259, I1372, I434, I1806, I2977, I1074, I4271, I4786, I50, I4009, I1476, I537, I3731, I1983, I2172, I4317, I2541, I163, I4970, I1737, I2805, I3322, I326, I2550, I4558, I2455, I2422, I1905, I1713, I4098, I3087, I1515, I1926, I2827, I4253, I1072, I2306, I3824, I2246, I506, I137, I3463, I2395, I2426, I1183, I4530, I123, I3244, I2751, I4596, I621, I816, I3124, I4475, I350, I4949, I4375, I2192, I15, I3219, I53, I2945, I3157, I2456, I619, I4774, I1558, I1606, I2158, I1274, I4025, I4026, I2864, I3599, I299, I583, I3497, I4164, I4086, I1493, I102, I2763, I1891, I3312, I2999, I420, I1047, I3419, I1206, I4612, I2024, I195, I3000, I1329, I4581, I3224, I1872, I1820, I3951, I1082, I1793, I512, I1432, I3620, I3355, I4213, I1555, I4144, I52, I149, I4006, I760, I3445, I3982, I4609, I4664, I2052, I2218, I1236, I943, I3373, I2617, I3830, I2119, I4106, I2874, I4355, I3962, I371, I1087, I1990, I462, I3144, I1184, I549, I4361, I1062, I2424, I4823, I4061, I1565, I4209, I540, I1698, I4647, I4722, I1744, I3790, I3495, I268, I4237, I724, I4228, I3403, I439, I505, I482, I3041, I894, I4892, I1632, I3950, I2412, I3776, I4081, I978, I4613, I4395, I2949, I223, I2199, I4700, I2983, I878, I1462, I1319, I1467, I1150, I3461, I1201, I4140, I4479, I2877, I460, I4396, I2664, I2733, I3747, I2755, I2338, I2255, I4497, I2575, I4402, I489, I3800, I3573, I4814, I38, I2992, I2055, I1063, I1007, I2123, I2556, I2568, I125, I2089, I1512, I1941, I4535, I4204, I182, I3546, I964, I97, I1984, I4073, I946, I2842, I3572, I4043, I1701, I1065, I4638, I4994, I4451, I2128, I1280, I4943, I1804, I2321, I2793, I4606, I4947, I3805, I3764, I1910, I4901, I1191, I3635, I178, I1377, I1037, I987, I3683, I1187, I222, I830, I3035, I1935, I3877, I2860, I374, I2916, I2332, I4280, I4968, I965, I4797, I3038, I2025, I1375, I1014, I831, I938, I2566, I1270, I3952, I2646, I2259, I1848, I2191, I4708, I4157, I2802, I4118, I199, I3979, I976, I4462, I805, I899, I4531, I3136, I3291, I1438, I3865, I1832, I3195, I4453, I4354, I2804, I625, I4501, I1874, I4373, I1244, I1854, I1695, I2066, I359, I1745, I2626, I1549, I2054, I1578, I3631, I2783, I2516, I1639, I150, I2728, I3352, I3342, I2640, I2790, I3208, I4150, I1653, I1754, I4608, I2535, I1262, I2553, I496, I4742, I2226, I687, I1895, I3002, I838, I3646, I4397, I2461, I1743, I1427, I680, I1002, I3405, I2240, I3205, I121, I4252, I892, I4168, I2271, I1894, I3271, I202, I1667, I726, I2281, I2393, I1302, I2439, I2413, I3821, I2001, I4363, I2245, I4064, I3006, I4302, I1612, I3767, I4393, I2644, I2667, I3526, I1696, I317, I2771, I2546, I1416, I269, I1989, I2832, I1762, I4749, I936, I3727, I4867, I963, I3159, I1442, I3099, I4791, I4339, I3841, I4663, I4362, I183, I1154, I1054, I2115, I3225, I2803, I4852, I738, I3390, I3453, I1028, I2153, I4940, I4747, I1547, I4292, I1449, I1672, I3344, I1490, I3274, I4429, I4955, I4100, I3524, I638, I1814, I2991, I2649, I1849, I416, I1221, I4903, I3993, I4218, I4572, I2331, I2583, I2170, I65, I1507, I4788, I3364, I693, I3826, I646, I2812, I1537, I72, I4040, I166, I2236, I1444, I3783, I116, I147, I1608, I3838, I3914, I3897, I763, I4678, I4019, I3912, I4967, I3003, I3210, I1138, I4338, I1657, I2387, I1009, I2839, I287, I377, I1234, I4262, I2981, I2189, I1686, I835, I3947, I2840, I1304, I3915, I4191, I4848, I2408, I4584, I4039, I459, I1031, I1480, I3744, I3652, I2539, I2197, I1139, I303, I3351, I516, I3241, I2750, I4246, I4551, I4411, I4022, I3109, I261, I2538, I545, I4084, I2122, I1883, I1341, I1101, I1587, I2307, I1254, I1550, I385, I3740, I1214, I2190, I1720, I574, I4463, I1534, I2656, I1589, I981, I3277, I2019, I4005, I3743, I813, I200, I649, I755, I2620, I473, I3801, I1396, I1220, I4662, I3012, I260, I4374, I2822, I3211, I3121, I298, I589, I32, I2410, I1772, I1010, I2986, I4953, I1760, I3926, I4320, I2434, I801, I562, I1734, I3890, I3226, I230, I3695, I2551, I3212, I1809, I1121, I4937, I4240, I592, I857, I2960, I2322, I564, I4560, I2509, I450, I4681, I3213, I1914, I1251, I4855, I3658, I1272, I1888, I3678, I2935, I1776, I1478, I1980, I2703, I563, I4137, I1598, I3350, I1094, I4036, I2282, I4723, I4817, I3261, I3730, I2665, I2660, I484, I747, I4784, I3794, I1584, I2091, I3549, I2791, I1356, I4543, I2243, I1040, I3167, I1128, I4683, I1354, I107, I657, I4650, I2020, I4125, I1471, I4909, I1348, I3207, I17, I4733, I3014, I245, I4935, I40, I3067, I2782, I3612, I2230, I1137, I3119, I3255, I4709, I2504, I4089, I2324, I3761, I3220, I4864, I2639, I4768, I2294, I2544, I2502, I4055, I1650, I1690, I2258, I4380, I4419, I143, I4178, I4254, I1845, I319, I723, I302, I727, I4293, I3018, I4820, I1788, I2007, I2841, I3150, I1800, I1739, I2411, I1621, I4103, I1649, I2746, I3083, I4288, I190, I3095, I1135, I1453, I2699, I4825, I99, I4672, I879, I700, I2452, I4923, I3385, I4882, I3332, I2357, I3990, I4477, I4132, I1182, I916, I2908, I3742, I4286, I1861, I4952, I4537, I1299, I4017, I3769, I2863, I3908, I3432, I4104, I1564, I758, I608, I2820, I1297, I1303, I4736, I3605, I4776, I2959, I2698, I1887, I1169, I3222, I660, I4951, I4620, I3441, I474, I1585, I1520, I3173, I4074, I3437, I1273, I4887, I1192, I538, I4794, I733, I1851, I768, I2377, I566, I4128, I971, I231, I2386, I1342, I4273, I1424, I1456, I2163, I3377, I3885, I105, I3729, I4388, I4829, I2021, I953, I3585, I2990, I3875, I2299, I173, I4975, I654, I787, I2598, I2047, I4790, I3507, I1924, I2762, I1673, I1554, I2308, I1530, I2941, I1603, I2678, I626, I2441, I4115, I4202, I1967, I2873, I3837, I1846, I207, I2466, I547, I4912, I2375, I1475, I3019, I880, I3016, I3691, I4918, I2599, I2291, I3485, I3846, I4772, I648, I1783, I4279, I1885, I501, I2384, I2996, I796, I467, I2532, I1501, I2000, I928, I3587, I3290, I2786, I1133, I2653, I4470, I4299, I2445, I2881, I1913, I2608, I1359, I348, I4908, I1938, I1000, I4408, I3519, I2168, I2854, I2286, I2469, I3269, I4685, I3145, I3072, I406, I699, I1136, I1766, I4366, I4263, I1993, I1725, I2887, I351, I4574, I1871, I1526, I2527, I3553, I2015, I4993, I2187, I2084, I3789, I689, I550, I3543, I3610, I2925, I3182, I799, I26, I844, I655, I2711, I3665, I2614, I866, I1142, I1961, I2870, I1570, I4275, I4508, I3833, I2144, I902, I1583, I1008, I188, I3102, I867, I1747, I153, I967, I4311, I1269, I307, I1532, I3302, I66, I205, I2149, I146, I777, I3848, I4383, I247, I596, I3959, I1919, I4247, I951, I1199, I3194, I1626, I1369, I4425, I2071, I4510, I2349, I1610, I1940, I3276, I926, I2694, I2559, I4309, I2672, I390, I2801, I2922, I4433, I3843, I3842, I3864, I2679, I3972, I769, I3624, I4063, I2313, I3901, I2843, I3664, I652, I278, I3112, I1001, I4186, I14, I3985, I4194, I675, I113, I1830, I3933, I1912, I4899, I4082, I734, I3597, I1186, I1655, I3063, I3680, I3862, I4436, I2513, I544, I101, I2253, I4622, I2451, I1819, I2359, I138, I1922, I3421, I3732, I2277, I2695, I4313, I2723, I2506, I1708, I2006, I1177, I2490, I361, I3410, I2096, I2890, I2443, I642, I4384, I3529, I3868, I4352, I3048, I3389, I2718, I701, I2486, I4215, I4456, I3275, I4010, I706, I3452, I2104, I4591, I3407, I2351, I3857, I255, I1085, I1164, I4440, I1897, I1529, I4488, I2968, I4642, I4087, I4303, I2062, I2825, I4801, I4826, I2232, I4434, I3751, I4480, I3592, I4851, I1712, I812, I4900, I4099, I162, I2545, I134, I2911, I1873, I1158, I1322, I4412, I3337, I3158, I3856, I4704, I910, I671, I2561, I2972, I3492, I3938, I44, I184, I3125, I1218, I3137, I2673, I1952, I2563, I2984, I3499, I3763, I1056, I643, I131, I4404, I3870, I39, I4268, I4793, I659, I959, I2449, I1705, I4707, I3552, I1370, I1305, I3234, I111, I2067, I383, I1841, I3239, I1147, I674, I1151, I2244, I1357, I737, I370, I4670, I535, I4752, I881, I1548, I1207, I1358, I3369, I1620, I4871, I4448, I4189, I1787, I1997, I3713, I2752, I2520, I465, I3623, I3439, I581, I2923, I1278, I2621, I1903, I1238, I3462, I429, I2248, I4861, I2756, I3675, I3021, I1115, I3114, I3273, I4245, I1215, I415, I1865, I1607, I1797, I4753, I923, I542, I1468, I1668, I1472, I2896, I398, I2017, I254, I4656, I2263, I975, I49, I1170, I2214, I1328, I3135, I1927, I4582, I4834, I1893, I4671, I2571, I2398, I4351, I1615, I2346, I3723, I1242, I1078, I4139, I3490, I2799, I158, I4415, I4141, I1852, I1828, I2645, I2710, I409, I449, I1934, I548, I4188, I10, I2247, I3250, I632, I1860, I3986, I1429, I611, I3528, I4605, I4654, I1261, I731, I3104, I3169, I1609, I4406, I1360, I4312, I2807, I907, I3882, I4865, I1850, I2897, I1023, I1189, I1756, I2489, I3075, I3714, I3853, I209, I979, I3252, I3217, I253, I4435, I204, I4946, I2630, I639, I1367, I1366, I3133, I304, I2997, I4525, I1243, I1084, I3174, I672, I2402, I3965, I3504, I2943, I322, I3974, I4990, I2034, I893, I2862, I1784, I927, I1855, I3633, I3113, I2875, I4457, I2902, I330, I344, I2037, I2209, I3093, I714, I2953, I3816, I3039, I4283, I4836, I2603, I2884, I3032, I4117, I308, I4680, I2405, I3187, I3542, I4181, I2205, I1387, I4472, I4385, I3363, I1437, I4489, I3166, I4878, I1266, I4368, I1836, I543, I2589, I2220, I4595, I1509, I1835, I1733, I1200, I3388, I2809, I1452, I3895, I1166, I3548, I1802, I771, I2610, I579, I3567, I2365, I3218, I4564, I4512, I3556, I851, I430, I3745, I216, I1670, I2038, I1228, I2717, I1921, I3251, I3245, I664, I4133, I4906, I2760, I300, I2491, I2319, I1433, I2041, I514, I4597, I1789, I601, I4819, I21, I293, I584, I2181, I4658, I4636, I4281, I4325, I2938, I4085, I4534, I2810, I4314, I647, I3921, I3987, I1483, I4816, I1525, I3466, I218, I259, I4227, I3795, I2880, I4077, I2284, I3883, I1729, I895, I541, I2463, I4600, I4212, I1291, I846, I3139, I4003, I3802, I1077, I4335, I3770, I393, I1948, I3257, I476, I2249, I1638, I4559, I4423, I4466, I3676, I3293, I1179, I3451, I2403, I1340, I4430, I2966, I187, I3886, I3701, I4276, I4577, I1964, I4399, I2347, I3013, I2939, I598, I2889, I4547, I3247, I1947, I3127, I2982, I1969, I1248, I2558, I3532, I4874, I1837, I1344, I3057, I1911, I4321, I3128, I4914, I3431, I4449, I3107, I3080, I3069, I1378, I962, I2382, I470, I1404, I849, I1294, I3586, I3309, I3070, I2135, I2882, I637, I2142, I413, I942, I4207, I1202, I1130, I3033, I4919, I3436, I1310, I140, I376, I73, I4894, I36, I4305, I174, I1813, I1498, I3590, I4889, I536, I1389, I4358, I2231, I2063, I2915, I1519, I591, I3028, I1027, I1688, I2963, I480, I4174, I114, I2124, I2704, I4414, I1884, I3233, I2495, I1036, I522, I335, I3007, I373, I4756, I94, I911, I2278, I3022, I1579, I746, I367, I3494, I1976, I1562, I337, I4105, I3978, I2816, I2268, I2159, I4196, I1647, I3596, I360, I3828, I3516, I2161, I3715, I4971, I2528, I1778, I3430, I3467, I4746, I4593, I2360, I1808, I3330, I3008, I531, I4603, I3082, I2304, I3206, I2060, I4939, I824, I1049, I4386, I1286, I1484, I1419, I4618, I1740, I2885, I2018, I2719, I1779, I311, I3787, I532, I4703, I823, I1678, I1351, I3229, I2940, I1535, I1227, I3091, I3184, I2355, I2654, I770, I4154, I454, I528, I1518, I2344, I1684, I1481, I1728, I807, I2297, I1300, I3278, I1560, I2336, I571, I2302, I4996, I4327, I1822, I2143, I3356, I1943, I3286, I717, I2975, I2289, I3401, I381, I2295, I4973, I277, I4401, I2797, I1971, I1510, I437, I719, I640, I762, I669, I688, I2229, I870, I3081, I3289, I141, I1385, I1625, I595, I3367, I2138, I920, I2442, I3566, I3446, I2579, I3925, I2511, I481, I2836, I2976, I4122, I1577, I1373, I945, I3448, I1954, I3954, I4341, I1235, I3418, I1968, I3117, I4758, I4495, I258, I1916, I4241, I3707, I4661, I4127, I889, I4604, I3999, I4235, I2637, I4720, I4726, I3728, I3074, I4539, I4180, I3086, I4686, I407, I4527, I773, I3474, I2330, I718, I917, I1687, I2987, I103, I827, I2195, I4792, I1795, I2648, I1767, I2448, I4519, I2194, I3045, I3958, I3394, I4592, I3246, I2379, I56, I2894, I1582, I748, I508, I2048, I994, I630, I776, I4697, I1195, I636, I1131, I4278, I3384, I2687, I4058, I2798, I33, I4153, I3670, I229, I3847, I3263, I4308, I833, I3387, I3283, I4954, I605, I749, I4627, I4474, I1981, I4034, I705, I4744, I941, I2708, I4832, I3940, I4831, I1962, I3176, I2098, I590, I4166, I1960, I4083, I3788, I4713, I2970, I4750, I3522, I1685, I4929, I3957, I3428, I4367, I4390, I3618, I217, I2132, I4029, I3024, I2651, I1486, I1287, I3544, I1944, I1092, I1314, I3298, I2926, I2814, I4740, I730, I2692, I4350, I357, I4257, I2126, I1724, I3347, I2689, I2577, I3305, I2508, I4877, I3997, I1152, I2595, I4921, I4872, I2173, I2533, I4810, I4617, I4491, I1504, I4136, I3582, I2715, I4337, I3887, I4598, I1956, I3941, I3191, I527, I4344, I1249, I2436, I3177, I4381, I1443, I2808, I142, I4239, I4731, I1497, I4516, I4206, I2773, I681, I3984, I1403, I2593, I4725, I2661, I4847, I2775, I4205, I2878, I2498, I2329, I3967, I1083, I3498, I826, I1624, I1171, I1466, I3980, I3335, I4376, I4307, I614, I3354, I3478, I988, I4216, I2432, I1661, I2111, I2969, I1918, I3859, I3381, I2406, I3357, I2196, I940, I1569, I4159, I4770, I3238, I1987, I410, I3655, I4020, I707, I4042, I729, I1346, I3092, I3752, I3482, I818, I4977, I2310, I3977, I2266, I2446, I4296, I3930, I375, I4893, I1174, I2298, I3196, I485, I475, I3383, I486, I4193, I2954, I3382, I68, I1012, I3768, I2256, I3307, I4231, I3686, I1020, I1250, I725, I3471, I2200, I2622, I2264, I280, I4732, I3515, I3476, I286, I3129, I850, O489, O205, O311, O373, O422, O149, O448, O399, O301, O387, O24, O104, O377, O183, O497, O342, O107, O265, O185, O408, O124, O343, O152, O58, O392, O5, O172, O46, O189, O20, O291, O132, O248, O485, O61, O371, O487, O211, O56, O98, O82, O67, O436, O77, O26, O420, O37, O349, O430, O391, O286, O155, O112, O25, O425, O129, O243, O486, O72, O170, O117, O464, O319, O309, O4, O66, O288, O43, O483, O22, O415, O249, O410, O251, O465, O74, O60, O402, O414, O105, O427, O115, O406, O348, O467, O353, O73, O16, O380, O178, O197, O407, O134, O498, O293, O220, O231, O259, O457, O450, O429, O473, O445, O401, O219, O492, O396, O157, O295, O133, O493, O332, O180, O51, O382, O224, O47, O97, O241, O423, O275, O122, O195, O250, O49, O323, O269, O163, O29, O225, O165, O394, O254, O109, O346, O266, O167, O359, O147, O417, O34, O64, O80, O318, O326, O228, O351, O199, O138, O91, O452, O35, O100, O186, O393, O110, O274, O52, O300, O490, O298, O459, O463, O294, O312, O310, O169, O33, O461, O182, O358, O85, O344, O495, O478, O83, O145, O469, O292, O247, O426, O270, O337, O451, O154, O162, O32, O271, O84, O302, O368, O336, O7, O374, O447, O160, O198, O384, O413, O89, O395, O338, O214, O379, O121, O453, O123, O131, O252, O38, O41, O184, O139, O352, O36, O237, O321, O366, O102, O201, O240, O78, O113, O491, O9, O263, O235, O404, O411, O92, O238, O264, O421, O143, O12, O283, O281, O466, O314, O30, O494, O94, O306, O62, O363, O153, O272, O213, O383, O324, O106, O330, O161, O13, O95, O236, O341, O419, O246, O127, O191, O365, O126, O328, O188, O223, O354, O70, O279, O268, O116, O474, O468, O111, O17, O287, O428, O403, O282, O230, O280, O76, O81, O156, O166, O193, O175, O242, O222, O217, O315, O385, O325, O320, O444, O260, O434, O284, O446, O424, O221, O90, O135, O28, O313, O480, O88, O435, O442, O206, O190, O44, O475, O239, O125, O140, O48, O488, O45, O150, O53, O484, O79, O386, O177, O6, O229, O181, O210, O479, O471, O119, O278, O14, O144, O477, O8, O173, O39, O390, O151, O0, O208, O54, O472, O262, O31, O375, O23, O400, O255, O244, O470, O245, O273, O355, O148, O317, O86, O409, O304, O65, O55, O389, O40, O357, O176, O87, O218, O108, O418, O308, O50, O289, O256, O59, O93, O179, O305, O345, O276, O367, O204, O455, O297, O10, O261, O412, O335, O171, O350, O378, O3, O462, O431, O458, O258, O192, O234, O136, O381, O130, O303, O440, O257, O356, O15, O339, O99, O267, O376, O296, O216, O398, O331, O75, O443, O460, O42, O334, O397, O194, O362, O158, O11, O159, O372, O439, O347, O146, O476, O164, O19, O364, O21, O290, O499, O369, O187, O215, O432, O57, O196, O202, O441, O212, O128, O71, O437, O361, O456, O277, O203, O482, O103, O416, O481, O209, O168, O226, O101, O118, O360, O388, O322, O141, O232, O285, O370, O2, O307, O340, O18, O63, O1, O333, O233, O120, O329, O142, O27, O496, O227, O316, O438, O68, O69, O253, O96, O449, O200, O174, O454, O327, O114, O433, O207, O137, O405, O299);
	input I4737, I4052, I3510, I389, I2768, I29, I1544, I1759, I1646, I4182, I4743, I4001, I2233, I397, I425, I1494, I2103, I2521, I1222, I491, I1594, I900, I4728, I3598, I1718, I3047, I2709, I4555, I4806, I2484, I193, I4557, I3044, I2462, I192, I2748, I4692, I1021, I16, I282, I1699, I3402, I3118, I2732, I3270, I2113, I76, I2613, I1430, I3071, I1076, I2564, I915, I1601, I391, I2780, I379, I1870, I334, I1769, I4135, I2866, I4047, I4323, I1347, I3300, I1930, I3395, I2693, I3699, I2725, I3560, I4190, I4657, I1631, I3694, I2002, I815, I4439, I3306, I1977, I4928, I523, I2073, I4846, I3473, I4290, I3949, I4983, I736, I4109, I604, I559, I2735, I3152, I3700, I3372, I832, I3570, I767, I4835, I2086, I1840, I2785, I2666, I3575, I721, I4665, I417, I69, I3588, I1052, I2624, I422, I875, I817, I500, I3534, I766, I67, I534, I1185, I4594, I3781, I3009, I2094, I1410, I989, I1257, I2065, I4359, I3100, I22, I3973, I1237, I328, I1662, I848, I3684, I1447, I2675, I1230, I2378, I392, I1738, I4152, I3989, I242, I778, I2389, I2022, I1561, I3968, I2097, I3098, I2004, I555, I1099, I2117, I4272, I1203, I2154, I4626, I4891, I4481, I4220, I600, I2811, I2343, I4568, I1876, I2418, I4035, I458, I1775, I3696, I3379, I4391, I3942, I1233, I4711, I925, I2059, I1563, I3892, I4287, I686, I4645, I12, I754, I3654, I526, I4102, I1665, I408, I1771, I2043, I1479, I677, I226, I154, I3540, I1551, I4076, I2514, I587, I4773, I800, I4575, I3688, I2492, I3773, I4549, I4824, I4795, I4628, I77, I568, I2125, I1816, I1355, I4260, I2376, I2581, I513, I2013, I339, I691, I2929, I1654, I271, I2582, I3440, I3791, I774, I3444, I1461, I1024, I2177, I4176, I3660, I1379, I4432, I1781, I346, I1323, I3459, I1117, I4934, I1317, I2480, I4904, I3151, I2409, I3380, I2758, I2118, I4145, I3464, I1256, I197, I3414, I2734, I808, I775, I1285, I2280, I1420, I1463, I3134, I1393, I1900, I4156, I3256, I1426, I739, I3442, I997, I2927, I1831, I3852, I4357, I57, I2353, I3358, I4171, I906, I3627, I1627, I119, I2036, I1815, I4049, I1482, I1079, I2744, I3809, I63, I635, I3648, I2070, I1574, I1155, I3638, I3235, I4378, I4048, I764, I4101, I3333, I1440, I4590, I2267, I3906, I4057, I3879, I2106, I2179, I914, I3900, I2241, I4334, I2061, I3512, I2447, I2095, I1637, I3361, I369, I521, I2683, I1097, I1301, I3172, I1597, I1659, I4160, I2777, I3480, I859, I58, I4023, I913, I3777, I3317, I2202, I2659, I3636, I4079, I493, I4195, I443, I678, I3110, I3750, I208, I599, I3966, I2437, I1992, I2152, I2828, I1877, I1540, I4883, I2033, I1160, I3324, I4763, I2702, I1617, I3673, I2713, I4255, I239, I1572, I2146, I1826, I4546, I4243, I948, I306, I3943, I3025, I1473, I1335, I2458, I4392, I2743, I3720, I4879, I821, I2865, I1522, I4856, I991, I2433, I3817, I1418, I2032, I1863, I74, I1966, I4944, I1116, I4054, I2160, I3722, I620, I418, I2137, I4394, I1140, I3345, I2475, I2224, I1896, I1260, I3215, I3065, I3058, I2988, I1553, I3077, I2364, I2769, I2450, I1204, I3138, I1868, I2868, I4573, I1320, I3237, I3656, I3602, I3326, I2588, I4234, I4369, I4646, I3406, I2642, I950, I3936, I1353, I1867, I1899, I4332, I4119, I2121, I3893, I3188, I1382, I1383, I3719, I623, I3170, I2162, I3164, I742, I1327, I2861, I1223, I1298, I4129, I2906, I2093, I4146, I4343, I1488, I1096, I4844, I969, I1330, I4830, I1710, I3316, I4804, I3026, I2392, I4469, I176, I918, I2858, I4405, I148, I3198, I240, I497, I2691, I856, I331, I1409, I3577, I3523, I2503, I510, I3457, I4760, I1112, I4571, I1108, I1915, I977, I585, I3780, I3296, I3815, I18, I5, I3297, I1190, I2937, I3663, I1265, I3017, I1004, I3771, I2217, I3054, I4285, I1492, I4649, I2049, I1073, I4601, I2633, I3685, I3181, I4624, I3935, I929, I2647, I4110, I2730, I905, I3806, I4616, I1683, I2368, I4225, I332, I1679, I720, I2677, I95, I90, I1857, I1487, I227, I1752, I19, I1425, I400, I575, I3192, I2188, I3066, I2427, I2425, I3216, I2003, I695, I1817, I4120, I2112, I1, I4261, I3969, I71, I553, I3996, I3325, I4370, I586, I3328, I3513, I1811, I4655, I1307, I3488, I1229, I3231, I3413, I1061, I3617, I3162, I3336, I2222, I4630, I3782, I499, I4203, I1321, I1660, I312, I3521, I2416, I2303, I1792, I2635, I3346, I155, I3376, I842, I4933, I3839, I3576, I3353, I698, I4526, I970, I3059, I4041, I4075, I2213, I2272, I2903, I4714, I4751, I4371, I3661, I3301, I433, I96, I2957, I3863, I477, I1159, I713, I1325, I1034, I1842, I2540, I3185, I4324, I4467, I70, I380, I610, I1132, I1694, I2193, I1465, I4602, I2109, I2099, I179, I243, I4447, I1178, I3946, I3896, I2216, I2127, I1514, I954, I1127, I3284, I4200, I4674, I3020, I4515, I4828, I2438, I3561, I214, I782, I1963, I2697, I3165, I4910, I2576, I2051, I858, I1768, I2688, I1936, I2225, I2523, I4545, I2789, I3396, I703, I1750, I2435, I471, I1029, I876, I4956, I3496, I2373, I1645, I4294, I1311, I267, I786, I2479, I2145, I228, I4621, I451, I1496, I1834, I4690, I206, I3472, I464, I4745, I2722, I980, I934, I2834, I3486, I1081, I1794, I1349, I4873, I2573, I2682, I4163, I78, I4331, I4045, I1384, I631, I868, I4902, I4963, I1648, I1879, I2044, I3934, I3708, I3425, I3903, I1415, I2305, I606, I2965, I2947, I196, I4169, I4942, I3200, I4524, I3793, I3668, I1669, I2676, I4158, I4787, I3349, I3417, I2251, I4863, I2180, I4142, I440, I1240, I3535, I2342, I2481, I59, I1143, I1974, I2219, I1859, I191, I897, I1247, I1451, I4778, I4868, I3386, I2223, I2601, I3869, I1677, I3153, I4679, I845, I829, I1017, I4382, I662, I1853, I676, I1972, I820, I3659, I3904, I1546, I4148, I447, I185, I313, I2765, I1839, I2348, I2312, I244, I2337, I4066, I1557, I3115, I3508, I2547, I2369, I603, I3147, I1692, I2815, I3778, I1345, I3236, I1386, I3178, I2358, I27, I2388, I3243, I1071, I382, I756, I87, I4821, I2108, I3429, I890, I4409, I1716, I3203, I4880, I1777, I4849, I1368, I1068, I1422, I3929, I3280, I349, I2083, I4799, I3323, I4980, I588, I2706, I3649, I4161, I2028, I4666, I365, I1477, I3040, I709, I4107, I1395, I479, I1552, I1957, I1709, I355, I803, I4730, I1605, I120, I990, I573, I2962, I921, I4346, I3878, I1953, I2453, I2580, I386, I4712, I2354, I2570, I4112, I4976, I4802, I4611, I2849, I1157, I3538, I3850, I3703, I51, I3202, I4710, I2895, I2796, I4012, I1293, I4221, I1003, I3201, I1455, I784, I4689, I2907, I4259, I2993, I1333, I4192, I2627, I4936, I2471, I177, I2830, I3584, I2585, I2641, I3171, I1567, I1517, I2631, I580, I115, I1770, I2363, I1556, I3279, I2140, I2669, I3272, I3639, I292, I3907, I735, I4991, I2824, I4913, I3594, I3503, I1991, I1761, I2994, I3796, I509, I241, I3415, I3435, I2211, I4958, I1723, I1043, I931, I4619, I152, I3299, I3046, I2417, I1790, I3759, I3601, I4410, I2075, I34, I54, I325, I4924, I1401, I1721, I2320, I1458, I939, I219, I2339, I750, I3334, I2421, I3108, I1988, I1469, I2276, I2428, I1365, I3772, I3365, I1454, I2512, I4486, I3391, I1039, I4808, I2201, I2087, I3183, I4859, I1032, I565, I4170, I4473, I2716, I3739, I4452, I3976, I1596, I2472, I1524, I3860, I4113, I3458, I1907, I1255, I3669, I3580, I3536, I1805, I4961, I622, I2609, I1188, I4300, I412, I1622, I3155, I1057, I7, I1405, I935, I2727, I2129, I1955, I968, I4459, I891, I641, I1516, I1388, I757, I715, I1727, I2749, I4062, I3479, I2525, I2754, I3314, I250, I4815, I4199, I8, I1786, I225, I4803, I3619, I124, I362, I2517, I2872, I569, I402, I3775, I618, I4845, I3304, I4987, I1528, I1909, I996, I855, I539, I1212, I494, I722, I4684, I4698, I4886, I1176, I4926, I3651, I4027, I912, I4599, I1197, I321, I2753, I4464, I1022, I4030, I1693, I1643, I3836, I4905, I780, I490, I2586, I1119, I4217, I4542, I3160, I2707, I3266, I2150, I4328, I4484, I3578, I2327, I1600, I3798, I3705, I984, I1196, I3094, I3339, I4927, I2394, I3123, I3606, I694, I3103, I1880, I3667, I822, I2237, I305, I903, I4201, I4028, I2157, I1030, I1241, I644, I4282, I3554, I4850, I1090, I1098, I1436, I1765, I1827, I4291, I2680, I3792, I295, I3456, I3455, I3840, I3449, I4676, I3611, I4785, I702, I4925, I2290, I118, I704, I1807, I3928, I1089, I1226, I1216, I4126, I828, I3029, I3811, I577, I3484, I272, I1838, I4986, I3310, I3672, I144, I2531, I4695, I4111, I3709, I3366, I3438, I2166, I1576, I1134, I4884, I3268, I3149, I661, I4015, I3991, I1999, I4615, I3374, I4185, I3820, I2460, I2257, I4985, I2701, I4607, I2473, I1446, I1141, I81, I2203, I4007, I3393, I4513, I2287, I2419, I3559, I1939, I2893, I1381, I4056, I275, I4860, I1829, I2920, I262, I1168, I4578, I4356, I4437, I2430, I3533, I1296, I3988, I765, I3671, I3910, I4984, I4982, I4092, I2714, I1798, I104, I3193, I4498, I431, I264, I291, I3079, I3564, I2837, I4000, I2040, I1731, I1923, I2597, I310, I4544, I3514, I2846, I3628, I1315, I399, I1045, I546, I3050, I411, I3221, I1932, I1352, I2165, I3282, I1856, I1075, I2314, I790, I4400, I372, I435, I1890, I2014, I1394, I1275, I1527, I1470, I2844, I4496, I4857, I2221, I3827, I4438, I2956, I3916, I2311, I3692, I4070, I3116, I4264, I2578, I4506, I3359, I1545, I974, I4805, I3757, I3468, I1067, I2739, I3209, I2829, I4068, I4069, I456, I3142, I602, I198, I4890, I290, I358, I4969, I4648, I2850, I1059, I2139, I3084, I3995, I2069, I3971, I1566, I1541, I3641, I1308, I1613, I578, I2919, I3812, I692, I3873, I1931, I315, I1326, I4222, I3360, I3315, I2562, I3001, I186, I461, I2301, I2340, I3506, I3052, I793, I4389, I4197, I2604, I288, I684, I3591, I2254, I663, I1933, I2658, I2720, I1390, I2784, I2657, I3061, I232, I48, I1306, I2831, I937, I1644, I2309, I4304, I888, I1614, I3545, I3717, I4297, I3765, I252, I4522, I13, I1148, I453, I2077, I1580, I4050, I478, I1642, I792, I1336, I2974, I4008, I3822, I3888, I3630, I3060, I4417, I4640, I728, I1700, I814, I4210, I1086, I1364, I238, I2493, I4764, I4653, I2068, I220, I3593, I2400, I3056, I567, I3992, I1400, I4771, I1942, I933, I2605, I4096, I1149, I1016, I4885, I2296, I1995, I2989, I1658, I2238, I3122, I1267, I1284, I1290, I4211, I3653, I690, I1742, I904, I1146, I1799, I4783, I2035, I2515, I3861, I343, I2482, I2380, I1785, I4431, I2352, I2005, I3608, I1575, I404, I3932, I165, I133, I256, I1421, I4011, I1123, I341, I1033, I4719, I3481, I960, I883, I2101, I1782, I2334, I3970, I1125, I2198, I167, I819, I2134, I4669, I2574, I3712, I518, I2971, I4822, I4471, I4660, I4322, I3062, I992, I1866, I1773, I3015, I2662, I3530, I2026, I1864, I3168, I854, I4420, I79, I1702, I2274, I2909, I3944, I4915, I64, I2606, I2857, I347, I4298, I1489, I3963, I4734, I3416, I4277, I2148, I2361, I345, I4336, I4033, I3662, I2478, I3981, I1434, I2596, I2779, I388, I2090, I4548, I2273, I3931, I4659, I2260, I572, I1506, I1485, I3180, I4177, I2483, I1371, I3163, I2817, I4078, I2835, I1847, I1937, I4407, I2924, I189, I4570, I1951, I4465, I1445, I3232, I711, I4629, I4931, I273, I4038, I871, I2381, I1595, I2391, I4143, I3629, I172, I92, I1439, I2345, I3565, I863, I732, I3568, I1173, I3408, I3832, I4532, I1103, I4319, I3621, I670, I314, I4869, I2042, I4091, I3214, I3248, I4090, I444, I432, I3704, I551, I2818, I3738, I25, I1889, I1500, I4635, I2900, I446, I336, I2102, I615, I4762, I3397, I983, I2175, I3625, I212, I956, I1640, I2133, I2184, I169, I4838, I4789, I2944, I2300, I3918, I3616, I1929, I1239, I1818, I4966, I2958, I2612, I1904, I3657, I1292, I4348, I2485, I1878, I2859, I741, I1536, I4114, I570, I1959, I3899, I4625, I761, I3724, I1970, I4269, I1869, I353, I4862, I257, I1862, I492, I2474, I4576, I1590, I795, I1823, I3961, I1664, I2788, I2724, I4306, I1350, I1641, I919, I4002, I4493, I1726, I2465, I650, I2250, I1996, I1219, I4579, I1402, I4800, I3876, I1391, I4016, I561, I2147, I1309, I3362, I1633, I1751, I3557, I3945, I743, I213, I1162, I455, I1753, I3953, I3491, I2856, I3341, I4807, I594, I3956, I3562, I2092, I3068, I503, I108, I2350, I4643, I2464, I1051, I2904, I41, I396, I483, I4031, I3392, I3294, I853, I4779, I2726, I23, I164, I2534, I139, I2397, I4131, I2404, I2046, I3154, I665, I4833, I957, I1011, I1908, I2072, I745, I520, I3891, I1107, I1289, I1533, I2420, I2731, I2151, I3027, I4067, I877, I697, I4748, I126, I4775, I3810, I1571, I3537, I4208, I3319, I3259, I1372, I434, I1806, I2977, I1074, I4271, I4786, I50, I4009, I1476, I537, I3731, I1983, I2172, I4317, I2541, I163, I4970, I1737, I2805, I3322, I326, I2550, I4558, I2455, I2422, I1905, I1713, I4098, I3087, I1515, I1926, I2827, I4253, I1072, I2306, I3824, I2246, I506, I137, I3463, I2395, I2426, I1183, I4530, I123, I3244, I2751, I4596, I621, I816, I3124, I4475, I350, I4949, I4375, I2192, I15, I3219, I53, I2945, I3157, I2456, I619, I4774, I1558, I1606, I2158, I1274, I4025, I4026, I2864, I3599, I299, I583, I3497, I4164, I4086, I1493, I102, I2763, I1891, I3312, I2999, I420, I1047, I3419, I1206, I4612, I2024, I195, I3000, I1329, I4581, I3224, I1872, I1820, I3951, I1082, I1793, I512, I1432, I3620, I3355, I4213, I1555, I4144, I52, I149, I4006, I760, I3445, I3982, I4609, I4664, I2052, I2218, I1236, I943, I3373, I2617, I3830, I2119, I4106, I2874, I4355, I3962, I371, I1087, I1990, I462, I3144, I1184, I549, I4361, I1062, I2424, I4823, I4061, I1565, I4209, I540, I1698, I4647, I4722, I1744, I3790, I3495, I268, I4237, I724, I4228, I3403, I439, I505, I482, I3041, I894, I4892, I1632, I3950, I2412, I3776, I4081, I978, I4613, I4395, I2949, I223, I2199, I4700, I2983, I878, I1462, I1319, I1467, I1150, I3461, I1201, I4140, I4479, I2877, I460, I4396, I2664, I2733, I3747, I2755, I2338, I2255, I4497, I2575, I4402, I489, I3800, I3573, I4814, I38, I2992, I2055, I1063, I1007, I2123, I2556, I2568, I125, I2089, I1512, I1941, I4535, I4204, I182, I3546, I964, I97, I1984, I4073, I946, I2842, I3572, I4043, I1701, I1065, I4638, I4994, I4451, I2128, I1280, I4943, I1804, I2321, I2793, I4606, I4947, I3805, I3764, I1910, I4901, I1191, I3635, I178, I1377, I1037, I987, I3683, I1187, I222, I830, I3035, I1935, I3877, I2860, I374, I2916, I2332, I4280, I4968, I965, I4797, I3038, I2025, I1375, I1014, I831, I938, I2566, I1270, I3952, I2646, I2259, I1848, I2191, I4708, I4157, I2802, I4118, I199, I3979, I976, I4462, I805, I899, I4531, I3136, I3291, I1438, I3865, I1832, I3195, I4453, I4354, I2804, I625, I4501, I1874, I4373, I1244, I1854, I1695, I2066, I359, I1745, I2626, I1549, I2054, I1578, I3631, I2783, I2516, I1639, I150, I2728, I3352, I3342, I2640, I2790, I3208, I4150, I1653, I1754, I4608, I2535, I1262, I2553, I496, I4742, I2226, I687, I1895, I3002, I838, I3646, I4397, I2461, I1743, I1427, I680, I1002, I3405, I2240, I3205, I121, I4252, I892, I4168, I2271, I1894, I3271, I202, I1667, I726, I2281, I2393, I1302, I2439, I2413, I3821, I2001, I4363, I2245, I4064, I3006, I4302, I1612, I3767, I4393, I2644, I2667, I3526, I1696, I317, I2771, I2546, I1416, I269, I1989, I2832, I1762, I4749, I936, I3727, I4867, I963, I3159, I1442, I3099, I4791, I4339, I3841, I4663, I4362, I183, I1154, I1054, I2115, I3225, I2803, I4852, I738, I3390, I3453, I1028, I2153, I4940, I4747, I1547, I4292, I1449, I1672, I3344, I1490, I3274, I4429, I4955, I4100, I3524, I638, I1814, I2991, I2649, I1849, I416, I1221, I4903, I3993, I4218, I4572, I2331, I2583, I2170, I65, I1507, I4788, I3364, I693, I3826, I646, I2812, I1537, I72, I4040, I166, I2236, I1444, I3783, I116, I147, I1608, I3838, I3914, I3897, I763, I4678, I4019, I3912, I4967, I3003, I3210, I1138, I4338, I1657, I2387, I1009, I2839, I287, I377, I1234, I4262, I2981, I2189, I1686, I835, I3947, I2840, I1304, I3915, I4191, I4848, I2408, I4584, I4039, I459, I1031, I1480, I3744, I3652, I2539, I2197, I1139, I303, I3351, I516, I3241, I2750, I4246, I4551, I4411, I4022, I3109, I261, I2538, I545, I4084, I2122, I1883, I1341, I1101, I1587, I2307, I1254, I1550, I385, I3740, I1214, I2190, I1720, I574, I4463, I1534, I2656, I1589, I981, I3277, I2019, I4005, I3743, I813, I200, I649, I755, I2620, I473, I3801, I1396, I1220, I4662, I3012, I260, I4374, I2822, I3211, I3121, I298, I589, I32, I2410, I1772, I1010, I2986, I4953, I1760, I3926, I4320, I2434, I801, I562, I1734, I3890, I3226, I230, I3695, I2551, I3212, I1809, I1121, I4937, I4240, I592, I857, I2960, I2322, I564, I4560, I2509, I450, I4681, I3213, I1914, I1251, I4855, I3658, I1272, I1888, I3678, I2935, I1776, I1478, I1980, I2703, I563, I4137, I1598, I3350, I1094, I4036, I2282, I4723, I4817, I3261, I3730, I2665, I2660, I484, I747, I4784, I3794, I1584, I2091, I3549, I2791, I1356, I4543, I2243, I1040, I3167, I1128, I4683, I1354, I107, I657, I4650, I2020, I4125, I1471, I4909, I1348, I3207, I17, I4733, I3014, I245, I4935, I40, I3067, I2782, I3612, I2230, I1137, I3119, I3255, I4709, I2504, I4089, I2324, I3761, I3220, I4864, I2639, I4768, I2294, I2544, I2502, I4055, I1650, I1690, I2258, I4380, I4419, I143, I4178, I4254, I1845, I319, I723, I302, I727, I4293, I3018, I4820, I1788, I2007, I2841, I3150, I1800, I1739, I2411, I1621, I4103, I1649, I2746, I3083, I4288, I190, I3095, I1135, I1453, I2699, I4825, I99, I4672, I879, I700, I2452, I4923, I3385, I4882, I3332, I2357, I3990, I4477, I4132, I1182, I916, I2908, I3742, I4286, I1861, I4952, I4537, I1299, I4017, I3769, I2863, I3908, I3432, I4104, I1564, I758, I608, I2820, I1297, I1303, I4736, I3605, I4776, I2959, I2698, I1887, I1169, I3222, I660, I4951, I4620, I3441, I474, I1585, I1520, I3173, I4074, I3437, I1273, I4887, I1192, I538, I4794, I733, I1851, I768, I2377, I566, I4128, I971, I231, I2386, I1342, I4273, I1424, I1456, I2163, I3377, I3885, I105, I3729, I4388, I4829, I2021, I953, I3585, I2990, I3875, I2299, I173, I4975, I654, I787, I2598, I2047, I4790, I3507, I1924, I2762, I1673, I1554, I2308, I1530, I2941, I1603, I2678, I626, I2441, I4115, I4202, I1967, I2873, I3837, I1846, I207, I2466, I547, I4912, I2375, I1475, I3019, I880, I3016, I3691, I4918, I2599, I2291, I3485, I3846, I4772, I648, I1783, I4279, I1885, I501, I2384, I2996, I796, I467, I2532, I1501, I2000, I928, I3587, I3290, I2786, I1133, I2653, I4470, I4299, I2445, I2881, I1913, I2608, I1359, I348, I4908, I1938, I1000, I4408, I3519, I2168, I2854, I2286, I2469, I3269, I4685, I3145, I3072, I406, I699, I1136, I1766, I4366, I4263, I1993, I1725, I2887, I351, I4574, I1871, I1526, I2527, I3553, I2015, I4993, I2187, I2084, I3789, I689, I550, I3543, I3610, I2925, I3182, I799, I26, I844, I655, I2711, I3665, I2614, I866, I1142, I1961, I2870, I1570, I4275, I4508, I3833, I2144, I902, I1583, I1008, I188, I3102, I867, I1747, I153, I967, I4311, I1269, I307, I1532, I3302, I66, I205, I2149, I146, I777, I3848, I4383, I247, I596, I3959, I1919, I4247, I951, I1199, I3194, I1626, I1369, I4425, I2071, I4510, I2349, I1610, I1940, I3276, I926, I2694, I2559, I4309, I2672, I390, I2801, I2922, I4433, I3843, I3842, I3864, I2679, I3972, I769, I3624, I4063, I2313, I3901, I2843, I3664, I652, I278, I3112, I1001, I4186, I14, I3985, I4194, I675, I113, I1830, I3933, I1912, I4899, I4082, I734, I3597, I1186, I1655, I3063, I3680, I3862, I4436, I2513, I544, I101, I2253, I4622, I2451, I1819, I2359, I138, I1922, I3421, I3732, I2277, I2695, I4313, I2723, I2506, I1708, I2006, I1177, I2490, I361, I3410, I2096, I2890, I2443, I642, I4384, I3529, I3868, I4352, I3048, I3389, I2718, I701, I2486, I4215, I4456, I3275, I4010, I706, I3452, I2104, I4591, I3407, I2351, I3857, I255, I1085, I1164, I4440, I1897, I1529, I4488, I2968, I4642, I4087, I4303, I2062, I2825, I4801, I4826, I2232, I4434, I3751, I4480, I3592, I4851, I1712, I812, I4900, I4099, I162, I2545, I134, I2911, I1873, I1158, I1322, I4412, I3337, I3158, I3856, I4704, I910, I671, I2561, I2972, I3492, I3938, I44, I184, I3125, I1218, I3137, I2673, I1952, I2563, I2984, I3499, I3763, I1056, I643, I131, I4404, I3870, I39, I4268, I4793, I659, I959, I2449, I1705, I4707, I3552, I1370, I1305, I3234, I111, I2067, I383, I1841, I3239, I1147, I674, I1151, I2244, I1357, I737, I370, I4670, I535, I4752, I881, I1548, I1207, I1358, I3369, I1620, I4871, I4448, I4189, I1787, I1997, I3713, I2752, I2520, I465, I3623, I3439, I581, I2923, I1278, I2621, I1903, I1238, I3462, I429, I2248, I4861, I2756, I3675, I3021, I1115, I3114, I3273, I4245, I1215, I415, I1865, I1607, I1797, I4753, I923, I542, I1468, I1668, I1472, I2896, I398, I2017, I254, I4656, I2263, I975, I49, I1170, I2214, I1328, I3135, I1927, I4582, I4834, I1893, I4671, I2571, I2398, I4351, I1615, I2346, I3723, I1242, I1078, I4139, I3490, I2799, I158, I4415, I4141, I1852, I1828, I2645, I2710, I409, I449, I1934, I548, I4188, I10, I2247, I3250, I632, I1860, I3986, I1429, I611, I3528, I4605, I4654, I1261, I731, I3104, I3169, I1609, I4406, I1360, I4312, I2807, I907, I3882, I4865, I1850, I2897, I1023, I1189, I1756, I2489, I3075, I3714, I3853, I209, I979, I3252, I3217, I253, I4435, I204, I4946, I2630, I639, I1367, I1366, I3133, I304, I2997, I4525, I1243, I1084, I3174, I672, I2402, I3965, I3504, I2943, I322, I3974, I4990, I2034, I893, I2862, I1784, I927, I1855, I3633, I3113, I2875, I4457, I2902, I330, I344, I2037, I2209, I3093, I714, I2953, I3816, I3039, I4283, I4836, I2603, I2884, I3032, I4117, I308, I4680, I2405, I3187, I3542, I4181, I2205, I1387, I4472, I4385, I3363, I1437, I4489, I3166, I4878, I1266, I4368, I1836, I543, I2589, I2220, I4595, I1509, I1835, I1733, I1200, I3388, I2809, I1452, I3895, I1166, I3548, I1802, I771, I2610, I579, I3567, I2365, I3218, I4564, I4512, I3556, I851, I430, I3745, I216, I1670, I2038, I1228, I2717, I1921, I3251, I3245, I664, I4133, I4906, I2760, I300, I2491, I2319, I1433, I2041, I514, I4597, I1789, I601, I4819, I21, I293, I584, I2181, I4658, I4636, I4281, I4325, I2938, I4085, I4534, I2810, I4314, I647, I3921, I3987, I1483, I4816, I1525, I3466, I218, I259, I4227, I3795, I2880, I4077, I2284, I3883, I1729, I895, I541, I2463, I4600, I4212, I1291, I846, I3139, I4003, I3802, I1077, I4335, I3770, I393, I1948, I3257, I476, I2249, I1638, I4559, I4423, I4466, I3676, I3293, I1179, I3451, I2403, I1340, I4430, I2966, I187, I3886, I3701, I4276, I4577, I1964, I4399, I2347, I3013, I2939, I598, I2889, I4547, I3247, I1947, I3127, I2982, I1969, I1248, I2558, I3532, I4874, I1837, I1344, I3057, I1911, I4321, I3128, I4914, I3431, I4449, I3107, I3080, I3069, I1378, I962, I2382, I470, I1404, I849, I1294, I3586, I3309, I3070, I2135, I2882, I637, I2142, I413, I942, I4207, I1202, I1130, I3033, I4919, I3436, I1310, I140, I376, I73, I4894, I36, I4305, I174, I1813, I1498, I3590, I4889, I536, I1389, I4358, I2231, I2063, I2915, I1519, I591, I3028, I1027, I1688, I2963, I480, I4174, I114, I2124, I2704, I4414, I1884, I3233, I2495, I1036, I522, I335, I3007, I373, I4756, I94, I911, I2278, I3022, I1579, I746, I367, I3494, I1976, I1562, I337, I4105, I3978, I2816, I2268, I2159, I4196, I1647, I3596, I360, I3828, I3516, I2161, I3715, I4971, I2528, I1778, I3430, I3467, I4746, I4593, I2360, I1808, I3330, I3008, I531, I4603, I3082, I2304, I3206, I2060, I4939, I824, I1049, I4386, I1286, I1484, I1419, I4618, I1740, I2885, I2018, I2719, I1779, I311, I3787, I532, I4703, I823, I1678, I1351, I3229, I2940, I1535, I1227, I3091, I3184, I2355, I2654, I770, I4154, I454, I528, I1518, I2344, I1684, I1481, I1728, I807, I2297, I1300, I3278, I1560, I2336, I571, I2302, I4996, I4327, I1822, I2143, I3356, I1943, I3286, I717, I2975, I2289, I3401, I381, I2295, I4973, I277, I4401, I2797, I1971, I1510, I437, I719, I640, I762, I669, I688, I2229, I870, I3081, I3289, I141, I1385, I1625, I595, I3367, I2138, I920, I2442, I3566, I3446, I2579, I3925, I2511, I481, I2836, I2976, I4122, I1577, I1373, I945, I3448, I1954, I3954, I4341, I1235, I3418, I1968, I3117, I4758, I4495, I258, I1916, I4241, I3707, I4661, I4127, I889, I4604, I3999, I4235, I2637, I4720, I4726, I3728, I3074, I4539, I4180, I3086, I4686, I407, I4527, I773, I3474, I2330, I718, I917, I1687, I2987, I103, I827, I2195, I4792, I1795, I2648, I1767, I2448, I4519, I2194, I3045, I3958, I3394, I4592, I3246, I2379, I56, I2894, I1582, I748, I508, I2048, I994, I630, I776, I4697, I1195, I636, I1131, I4278, I3384, I2687, I4058, I2798, I33, I4153, I3670, I229, I3847, I3263, I4308, I833, I3387, I3283, I4954, I605, I749, I4627, I4474, I1981, I4034, I705, I4744, I941, I2708, I4832, I3940, I4831, I1962, I3176, I2098, I590, I4166, I1960, I4083, I3788, I4713, I2970, I4750, I3522, I1685, I4929, I3957, I3428, I4367, I4390, I3618, I217, I2132, I4029, I3024, I2651, I1486, I1287, I3544, I1944, I1092, I1314, I3298, I2926, I2814, I4740, I730, I2692, I4350, I357, I4257, I2126, I1724, I3347, I2689, I2577, I3305, I2508, I4877, I3997, I1152, I2595, I4921, I4872, I2173, I2533, I4810, I4617, I4491, I1504, I4136, I3582, I2715, I4337, I3887, I4598, I1956, I3941, I3191, I527, I4344, I1249, I2436, I3177, I4381, I1443, I2808, I142, I4239, I4731, I1497, I4516, I4206, I2773, I681, I3984, I1403, I2593, I4725, I2661, I4847, I2775, I4205, I2878, I2498, I2329, I3967, I1083, I3498, I826, I1624, I1171, I1466, I3980, I3335, I4376, I4307, I614, I3354, I3478, I988, I4216, I2432, I1661, I2111, I2969, I1918, I3859, I3381, I2406, I3357, I2196, I940, I1569, I4159, I4770, I3238, I1987, I410, I3655, I4020, I707, I4042, I729, I1346, I3092, I3752, I3482, I818, I4977, I2310, I3977, I2266, I2446, I4296, I3930, I375, I4893, I1174, I2298, I3196, I485, I475, I3383, I486, I4193, I2954, I3382, I68, I1012, I3768, I2256, I3307, I4231, I3686, I1020, I1250, I725, I3471, I2200, I2622, I2264, I280, I4732, I3515, I3476, I286, I3129, I850;
	output O489, O205, O311, O373, O422, O149, O448, O399, O301, O387, O24, O104, O377, O183, O497, O342, O107, O265, O185, O408, O124, O343, O152, O58, O392, O5, O172, O46, O189, O20, O291, O132, O248, O485, O61, O371, O487, O211, O56, O98, O82, O67, O436, O77, O26, O420, O37, O349, O430, O391, O286, O155, O112, O25, O425, O129, O243, O486, O72, O170, O117, O464, O319, O309, O4, O66, O288, O43, O483, O22, O415, O249, O410, O251, O465, O74, O60, O402, O414, O105, O427, O115, O406, O348, O467, O353, O73, O16, O380, O178, O197, O407, O134, O498, O293, O220, O231, O259, O457, O450, O429, O473, O445, O401, O219, O492, O396, O157, O295, O133, O493, O332, O180, O51, O382, O224, O47, O97, O241, O423, O275, O122, O195, O250, O49, O323, O269, O163, O29, O225, O165, O394, O254, O109, O346, O266, O167, O359, O147, O417, O34, O64, O80, O318, O326, O228, O351, O199, O138, O91, O452, O35, O100, O186, O393, O110, O274, O52, O300, O490, O298, O459, O463, O294, O312, O310, O169, O33, O461, O182, O358, O85, O344, O495, O478, O83, O145, O469, O292, O247, O426, O270, O337, O451, O154, O162, O32, O271, O84, O302, O368, O336, O7, O374, O447, O160, O198, O384, O413, O89, O395, O338, O214, O379, O121, O453, O123, O131, O252, O38, O41, O184, O139, O352, O36, O237, O321, O366, O102, O201, O240, O78, O113, O491, O9, O263, O235, O404, O411, O92, O238, O264, O421, O143, O12, O283, O281, O466, O314, O30, O494, O94, O306, O62, O363, O153, O272, O213, O383, O324, O106, O330, O161, O13, O95, O236, O341, O419, O246, O127, O191, O365, O126, O328, O188, O223, O354, O70, O279, O268, O116, O474, O468, O111, O17, O287, O428, O403, O282, O230, O280, O76, O81, O156, O166, O193, O175, O242, O222, O217, O315, O385, O325, O320, O444, O260, O434, O284, O446, O424, O221, O90, O135, O28, O313, O480, O88, O435, O442, O206, O190, O44, O475, O239, O125, O140, O48, O488, O45, O150, O53, O484, O79, O386, O177, O6, O229, O181, O210, O479, O471, O119, O278, O14, O144, O477, O8, O173, O39, O390, O151, O0, O208, O54, O472, O262, O31, O375, O23, O400, O255, O244, O470, O245, O273, O355, O148, O317, O86, O409, O304, O65, O55, O389, O40, O357, O176, O87, O218, O108, O418, O308, O50, O289, O256, O59, O93, O179, O305, O345, O276, O367, O204, O455, O297, O10, O261, O412, O335, O171, O350, O378, O3, O462, O431, O458, O258, O192, O234, O136, O381, O130, O303, O440, O257, O356, O15, O339, O99, O267, O376, O296, O216, O398, O331, O75, O443, O460, O42, O334, O397, O194, O362, O158, O11, O159, O372, O439, O347, O146, O476, O164, O19, O364, O21, O290, O499, O369, O187, O215, O432, O57, O196, O202, O441, O212, O128, O71, O437, O361, O456, O277, O203, O482, O103, O416, O481, O209, O168, O226, O101, O118, O360, O388, O322, O141, O232, O285, O370, O2, O307, O340, O18, O63, O1, O333, O233, O120, O329, O142, O27, O496, O227, O316, O438, O68, O69, O253, O96, O449, O200, O174, O454, O327, O114, O433, O207, O137, O405, O299;
	wire W0, W2, W5, W8, W9, W10, W11, W12, W17, W18, W21, W22, W25, W33, W35, W36, W39, W40, W41, W45, W47, W50, W53, W57, W58, W63, W68, W69, W72, W73, W74, W85, W88, W90, W91, W92, W94, W96, W98, W102, W106, W107, W108, W112, W113, W114, W117, W119, W120, W121, W122, W125, W126, W127, W129, W132, W136, W137, W138, W140, W144, W150, W151, W152, W153, W155, W156, W157, W159, W161, W162, W166, W175, W176, W180, W185, W188, W189, W191, W193, W195, W196, W198, W199, W201, W204, W205, W207, W212, W215, W217, W220, W223, W224, W229, W236, W246, W248, W249, W256, W260, W264, W265, W273, W276, W277, W278, W284, W285, W289, W297, W303, W304, W305, W306, W311, W318, W319, W322, W323, W324, W325, W327, W330, W336, W341, W344, W345, W347, W352, W355, W357, W358, W360, W370, W374, W378, W382, W388, W391, W394, W398, W400, W404, W405, W408, W409, W411, W414, W418, W419, W423, W424, W426, W428, W430, W432, W433, W437, W440, W441, W442, W445, W446, W447, W449, W450, W451, W453, W456, W458, W459, W463, W466, W468, W470, W471, W476, W479, W481, W486, W487, W488, W493, W497, W498, W499, W504, W510, W513, W515, W516, W517, W519, W526, W528, W529, W531, W533, W534, W536, W537, W541, W547, W548, W556, W564, W565, W568, W571, W575, W577, W581, W582, W585, W589, W593, W595, W596, W599, W600, W603, W604, W606, W607, W614, W617, W619, W621, W624, W625, W626, W630, W631, W633, W634, W635, W637, W638, W639, W640, W642, W646, W649, W652, W660, W661, W664, W665, W667, W671, W674, W676, W683, W686, W691, W693, W697, W702, W707, W711, W712, W713, W716, W720, W728, W729, W731, W735, W745, W747, W748, W750, W756, W757, W759, W760, W764, W766, W771, W775, W776, W782, W783, W784, W785, W786, W787, W788, W791, W792, W796, W797, W800, W802, W803, W805, W807, W811, W826, W831, W833, W837, W838, W840, W841, W842, W848, W854, W856, W860, W864, W869, W873, W878, W879, W881, W882, W884, W885, W888, W890, W896, W898, W899, W901, W902, W904, W908, W909, W913, W914, W915, W918, W924, W926, W929, W932, W935, W942, W944, W952, W954, W957, W959, W960, W964, W972, W973, W976, W977, W980, W982, W983, W984, W985, W987, W988, W991, W992, W1002, W1004, W1012, W1014, W1016, W1019, W1026, W1027, W1028, W1033, W1036, W1037, W1038, W1039, W1040, W1044, W1045, W1048, W1050, W1059, W1061, W1064, W1065, W1066, W1067, W1069, W1079, W1085, W1091, W1092, W1095, W1096, W1097, W1108, W1113, W1117, W1118, W1120, W1126, W1133, W1138, W1139, W1140, W1145, W1153, W1154, W1158, W1160, W1168, W1172, W1178, W1179, W1182, W1185, W1186, W1188, W1189, W1190, W1192, W1194, W1201, W1205, W1211, W1214, W1216, W1218, W1219, W1225, W1231, W1233, W1234, W1237, W1241, W1242, W1247, W1251, W1253, W1272, W1273, W1274, W1275, W1284, W1285, W1289, W1291, W1292, W1293, W1297, W1301, W1304, W1311, W1319, W1320, W1322, W1324, W1326, W1328, W1329, W1334, W1339, W1341, W1344, W1345, W1351, W1353, W1357, W1363, W1370, W1372, W1373, W1374, W1377, W1380, W1381, W1382, W1386, W1387, W1388, W1389, W1392, W1396, W1399, W1400, W1401, W1405, W1408, W1410, W1411, W1415, W1416, W1417, W1420, W1425, W1430, W1433, W1434, W1439, W1454, W1458, W1462, W1469, W1470, W1473, W1474, W1476, W1477, W1482, W1489, W1490, W1495, W1496, W1502, W1503, W1509, W1517, W1519, W1523, W1527, W1528, W1536, W1537, W1538, W1539, W1540, W1541, W1548, W1558, W1561, W1562, W1564, W1566, W1567, W1568, W1571, W1574, W1581, W1585, W1589, W1592, W1593, W1598, W1604, W1610, W1620, W1624, W1633, W1637, W1642, W1655, W1656, W1657, W1659, W1661, W1672, W1673, W1679, W1680, W1688, W1690, W1691, W1693, W1697, W1698, W1714, W1718, W1719, W1720, W1721, W1725, W1726, W1732, W1736, W1737, W1741, W1742, W1744, W1747, W1761, W1762, W1763, W1767, W1769, W1770, W1772, W1774, W1779, W1781, W1785, W1795, W1797, W1799, W1801, W1802, W1813, W1815, W1821, W1823, W1834, W1837, W1844, W1850, W1863, W1864, W1868, W1874, W1881, W1886, W1890, W1895, W1910, W1913, W1915, W1918, W1923, W1927, W1930, W1931, W1932, W1934, W1942, W1944, W1946, W1948, W1951, W1956, W1959, W1960, W1961, W1963, W1966, W1970, W1976, W1980, W1981, W1982, W1998, W2005, W2007, W2010, W2012, W2018, W2019, W2031, W2035, W2040, W2045, W2047, W2048, W2050, W2053, W2057, W2061, W2066, W2070, W2072, W2080, W2083, W2085, W2087, W2093, W2099, W2101, W2103, W2115, W2121, W2131, W2136, W2138, W2142, W2144, W2146, W2147, W2151, W2154, W2169, W2171, W2178, W2183, W2184, W2188, W2189, W2194, W2196, W2203, W2208, W2212, W2216, W2223, W2225, W2230, W2235, W2237, W2239, W2247, W2254, W2259, W2264, W2266, W2267, W2277, W2278, W2282, W2283, W2293, W2294, W2296, W2297, W2298, W2302, W2313, W2316, W2320, W2321, W2327, W2329, W2331, W2335, W2339, W2340, W2341, W2343, W2346, W2349, W2354, W2362, W2375, W2382, W2386, W2387, W2389, W2392, W2394, W2398, W2400, W2403, W2408, W2410, W2411, W2413, W2416, W2418, W2422, W2427, W2436, W2438, W2439, W2441, W2453, W2455, W2456, W2465, W2468, W2472, W2476, W2480, W2483, W2487, W2488, W2489, W2493, W2497, W2498, W2507, W2513, W2514, W2525, W2528, W2547, W2552, W2555, W2561, W2573, W2577, W2579, W2584, W2587, W2589, W2598, W2604, W2620, W2622, W2627, W2628, W2630, W2634, W2637, W2648, W2650, W2653, W2668, W2670, W2671, W2676, W2682, W2683, W2689, W2690, W2691, W2692, W2696, W2697, W2713, W2718, W2723, W2725, W2727, W2745, W2753, W2754, W2757, W2758, W2764, W2771, W2775, W2783, W2786, W2789, W2792, W2798, W2803, W2806, W2818, W2828, W2831, W2835, W2837, W2842, W2864, W2881, W2889, W2903, W2910, W2928, W2933, W2937, W2955, W2957, W2958, W2964, W2973, W2974, W2979, W2984, W2987, W3002, W3005, W3013, W3014, W3021, W3023, W3032, W3036, W3037, W3052, W3053, W3066, W3072, W3075, W3083, W3084, W3089, W3090, W3099, W3104, W3105, W3110, W3126, W3127, W3132, W3137, W3138, W3141, W3144, W3159, W3164, W3176, W3185, W3192, W3203, W3205, W3215, W3216, W3226, W3227, W3229, W3237, W3246, W3247, W3250, W3261, W3265, W3271, W3278, W3282, W3288, W3289, W3298, W3301, W3302, W3317, W3318, W3333, W3344, W3352, W3363, W3368, W3376, W3380, W3381, W3400, W3405, W3430, W3435, W3441, W3445, W3448, W3449, W3450, W3452, W3453, W3457, W3464, W3481, W3495, W3497, W3502, W3520, W3535, W3560, W3562, W3565, W3566, W3572, W3584, W3591, W3627, W3629, W3632, W3636, W3637, W3639, W3645, W3646, W3647, W3657, W3659, W3663, W3664, W3667, W3677, W3686, W3698, W3699, W3704, W3712, W3717, W3718, W3723, W3734, W3790, W3799, W3809, W3810, W3815, W3816, W3827, W3833, W3842, W3843, W3847, W3849, W3852, W3859, W3860, W3867, W3868, W3873, W3878, W3897, W3913, W3923, W3924, W3928, W3937, W3939, W3942, W3950, W3953, W3955, W3968, W3970, W3974, W3983, W3986, W3991, W3993, W3994, W3999, W4004, W4017, W4033, W4035, W4063, W4065, W4079, W4083, W4084, W4097, W4112, W4113, W4115, W4118, W4121, W4129, W4131, W4138, W4139, W4163, W4164, W4214, W4229, W4259, W4264, W4267, W4271, W4283, W4294, W4296, W4302, W4304, W4305, W4323, W4325, W4334, W4347, W4357, W4367, W4412, W4414, W4421, W4423, W4433, W4435, W4438, W4440, W4451, W4453, W4466, W4468, W4476, W4478, W4488, W4499, W4508, W4516, W4517, W4552, W4572, W4573, W4597, W4598, W4601, W4607, W4608, W4619, W4626, W4630, W4635, W4638, W4651, W4657, W4673, W4688, W4697, W4706, W4738, W4754, W4794, W4799, W4822, W4824, W4828, W4831, W4865, W4883, W4886, W4909, W4919, W4920, W4938, W4947, W4959, W4962, W4965, W4966, W4985, W4991, W4993, W5009, W5013, W5027, W5036, W5049, W5054, W5069, W5073, W5088, W5099, W5101, W5113, W5117, W5125, W5153, W5174, W5197, W5211, W5229, W5231, W5233, W5235, W5241, W5276, W5278, W5283, W5324, W5327, W5333, W5334, W5336, W5356, W5363, W5372, W5373, W5375, W5378, W5382, W5388, W5403, W5404, W5405, W5426, W5427, W5437, W5467, W5487, W5513, W5515, W5533, W5546, W5559, W5587, W5618, W5664, W5683, W5709, W5715, W5730, W5743, W5790, W5799, W5827, W5846, W5886, W5911, W5922, W5951, W5953, W5959, W5978, W5982, W5989, W5996, W5999, W6035, W6053, W6083, W6086, W6087, W6100, W6118, W6145, W6173, W6204, W6262, W6278, W6292, W6314, W6320, W6375, W6382, W6383, W6386, W6391, W6403, W6406, W6408, W6417, W6431, W6455, W6476, W6512, W6524, W6533, W6559, W6572, W6586, W6594, W6636, W6740, W6746, W6765, W6782, W6801, W6807, W6820, W6824, W6875, W6902, W6953, W6957, W6987, W6988, W7023, W7042, W7127, W7145, W7154, W7241, W7347, W7351, W7377, W7381, W7433, W7446, W7463, W7519, W7529, W7592, W7678, W7752, W7880, W7917, W7959, W8008, W8095, W8167, W8231, W8351, W8476, W8485, W8506, W8635, W8795, W9118, W9134, W9213;

	NANDX1 U0 (.A1(I3675), .A2(I967), .ZN(W0));
	NOR2X1 U2 (.A1(I1206), .A2(I1899), .ZN(W2));
	NOR2X1 U5 (.A1(I992), .A2(I1778), .ZN(W5));
	NOR2X1 U7 (.A1(I1695), .A2(I2982), .ZN(O44));
	NOR2X1 U8 (.A1(I801), .A2(I4908), .ZN(W8));
	NOR2X1 U9 (.A1(I4464), .A2(I3712), .ZN(W9));
	NOR2X1 U10 (.A1(I3723), .A2(I4156), .ZN(W10));
	INVX1 U11 (.I(I3087), .ZN(W11));
	INVX1 U12 (.I(I1525), .ZN(W12));
	NOR2X1 U13 (.A1(I252), .A2(I1536), .ZN(O330));
	NOR2X1 U17 (.A1(I1960), .A2(I1234), .ZN(W17));
	NANDX1 U18 (.A1(I4085), .A2(I1512), .ZN(W18));
	INVX1 U21 (.I(I4139), .ZN(W21));
	NOR2X1 U22 (.A1(I2647), .A2(I2963), .ZN(W22));
	NOR2X1 U25 (.A1(I1836), .A2(I2104), .ZN(W25));
	NANDX1 U33 (.A1(I176), .A2(I4350), .ZN(W33));
	NOR2X1 U35 (.A1(I3225), .A2(I823), .ZN(W35));
	NANDX1 U36 (.A1(I2990), .A2(I2284), .ZN(W36));
	NANDX1 U38 (.A1(I2958), .A2(I2005), .ZN(O408));
	INVX1 U39 (.I(I2656), .ZN(W39));
	NANDX1 U40 (.A1(I2699), .A2(I2640), .ZN(W40));
	NANDX1 U41 (.A1(I3436), .A2(I409), .ZN(W41));
	NANDX1 U45 (.A1(I1798), .A2(I3446), .ZN(W45));
	NOR2X1 U47 (.A1(I939), .A2(I4337), .ZN(W47));
	INVX1 U50 (.I(I4872), .ZN(W50));
	NOR2X1 U53 (.A1(I1836), .A2(I355), .ZN(W53));
	NANDX1 U57 (.A1(I2128), .A2(I3174), .ZN(W57));
	NOR2X1 U58 (.A1(I3316), .A2(I1135), .ZN(W58));
	NOR2X1 U63 (.A1(I4658), .A2(I1470), .ZN(W63));
	NOR2X1 U68 (.A1(I3169), .A2(I1395), .ZN(W68));
	NANDX1 U69 (.A1(I41), .A2(I1037), .ZN(W69));
	INVX1 U70 (.I(I4750), .ZN(O381));
	NOR2X1 U72 (.A1(I1778), .A2(I4770), .ZN(W72));
	NANDX1 U73 (.A1(I4477), .A2(I2662), .ZN(W73));
	NOR2X1 U74 (.A1(I3940), .A2(I1934), .ZN(W74));
	NANDX1 U85 (.A1(I4357), .A2(I3770), .ZN(W85));
	INVX1 U88 (.I(I968), .ZN(W88));
	NANDX1 U90 (.A1(I1421), .A2(I111), .ZN(W90));
	NANDX1 U91 (.A1(I1790), .A2(I4709), .ZN(W91));
	NANDX1 U92 (.A1(I1149), .A2(I3883), .ZN(W92));
	NOR2X1 U94 (.A1(I2972), .A2(I3655), .ZN(W94));
	NANDX1 U96 (.A1(I3191), .A2(I4041), .ZN(W96));
	INVX1 U98 (.I(I1553), .ZN(W98));
	NANDX1 U102 (.A1(I583), .A2(I4859), .ZN(W102));
	NANDX1 U106 (.A1(I2273), .A2(I2452), .ZN(W106));
	NANDX1 U107 (.A1(I3982), .A2(I535), .ZN(W107));
	NOR2X1 U108 (.A1(I1158), .A2(I1192), .ZN(W108));
	NOR2X1 U111 (.A1(W41), .A2(I3457), .ZN(O482));
	NOR2X1 U112 (.A1(I4513), .A2(I1626), .ZN(W112));
	NOR2X1 U113 (.A1(I835), .A2(I3883), .ZN(W113));
	NANDX1 U114 (.A1(I2953), .A2(I450), .ZN(W114));
	NANDX1 U117 (.A1(I3003), .A2(I2896), .ZN(W117));
	INVX1 U119 (.I(I3795), .ZN(W119));
	NANDX1 U120 (.A1(I991), .A2(I4790), .ZN(W120));
	INVX1 U121 (.I(I2775), .ZN(W121));
	NOR2X1 U122 (.A1(I725), .A2(I3133), .ZN(W122));
	INVX1 U125 (.I(I2249), .ZN(W125));
	NOR2X1 U126 (.A1(I4508), .A2(I1489), .ZN(W126));
	NOR2X1 U127 (.A1(I1401), .A2(I4579), .ZN(W127));
	NOR2X1 U129 (.A1(I3128), .A2(I462), .ZN(W129));
	NOR2X1 U130 (.A1(I941), .A2(I1747), .ZN(O487));
	NOR2X1 U132 (.A1(I1888), .A2(I4789), .ZN(W132));
	NOR2X1 U136 (.A1(I2035), .A2(I2831), .ZN(W136));
	NANDX1 U137 (.A1(I2268), .A2(I1923), .ZN(W137));
	NOR2X1 U138 (.A1(I799), .A2(I4661), .ZN(W138));
	NOR2X1 U140 (.A1(I335), .A2(I4111), .ZN(W140));
	NANDX1 U144 (.A1(I827), .A2(I3680), .ZN(W144));
	NOR2X1 U150 (.A1(I1486), .A2(I3294), .ZN(W150));
	NANDX1 U151 (.A1(I569), .A2(I3545), .ZN(W151));
	NOR2X1 U152 (.A1(I1900), .A2(I4040), .ZN(W152));
	NOR2X1 U153 (.A1(I1485), .A2(I1756), .ZN(W153));
	NOR2X1 U155 (.A1(I671), .A2(I4381), .ZN(W155));
	INVX1 U156 (.I(I1228), .ZN(W156));
	INVX1 U157 (.I(W68), .ZN(W157));
	NOR2X1 U159 (.A1(I1819), .A2(I3002), .ZN(W159));
	INVX1 U161 (.I(I4816), .ZN(W161));
	NANDX1 U162 (.A1(I793), .A2(I3128), .ZN(W162));
	NANDX1 U165 (.A1(I2392), .A2(I2935), .ZN(O72));
	INVX1 U166 (.I(I166), .ZN(W166));
	NANDX1 U174 (.A1(I1625), .A2(I3304), .ZN(O136));
	NOR2X1 U175 (.A1(I1738), .A2(I1787), .ZN(W175));
	NOR2X1 U176 (.A1(I4993), .A2(I4990), .ZN(W176));
	NOR2X1 U180 (.A1(I310), .A2(I564), .ZN(W180));
	NOR2X1 U185 (.A1(I2960), .A2(I4425), .ZN(W185));
	INVX1 U188 (.I(W132), .ZN(W188));
	NOR2X1 U189 (.A1(I4784), .A2(I95), .ZN(W189));
	INVX1 U191 (.I(I551), .ZN(W191));
	NOR2X1 U193 (.A1(I1809), .A2(I807), .ZN(W193));
	NANDX1 U195 (.A1(I747), .A2(I2231), .ZN(W195));
	NANDX1 U196 (.A1(I437), .A2(I4154), .ZN(W196));
	NANDX1 U198 (.A1(I3568), .A2(I1221), .ZN(W198));
	NANDX1 U199 (.A1(I123), .A2(I4534), .ZN(W199));
	INVX1 U201 (.I(I4158), .ZN(W201));
	NOR2X1 U204 (.A1(I505), .A2(I2754), .ZN(W204));
	NOR2X1 U205 (.A1(I2857), .A2(I4884), .ZN(W205));
	NANDX1 U207 (.A1(I1924), .A2(I3544), .ZN(W207));
	NOR2X1 U212 (.A1(I4117), .A2(I1270), .ZN(W212));
	NANDX1 U215 (.A1(I1151), .A2(I490), .ZN(W215));
	NANDX1 U217 (.A1(I485), .A2(I3008), .ZN(W217));
	NANDX1 U220 (.A1(I723), .A2(W175), .ZN(W220));
	NANDX1 U221 (.A1(I3451), .A2(I1150), .ZN(O296));
	INVX1 U223 (.I(I3229), .ZN(W223));
	NANDX1 U224 (.A1(I231), .A2(I631), .ZN(W224));
	INVX1 U229 (.I(I3620), .ZN(W229));
	NOR2X1 U236 (.A1(I1776), .A2(I1872), .ZN(W236));
	INVX1 U237 (.I(I3357), .ZN(O77));
	NANDX1 U242 (.A1(I3792), .A2(I2990), .ZN(O75));
	NOR2X1 U246 (.A1(I1911), .A2(I454), .ZN(W246));
	NANDX1 U248 (.A1(I2627), .A2(I169), .ZN(W248));
	INVX1 U249 (.I(I1496), .ZN(W249));
	INVX1 U252 (.I(I824), .ZN(O88));
	NOR2X1 U256 (.A1(I4596), .A2(W236), .ZN(W256));
	INVX1 U260 (.I(I4712), .ZN(W260));
	INVX1 U264 (.I(I877), .ZN(W264));
	NANDX1 U265 (.A1(W191), .A2(I2920), .ZN(W265));
	NOR2X1 U273 (.A1(W136), .A2(I3478), .ZN(W273));
	INVX1 U276 (.I(I174), .ZN(W276));
	NOR2X1 U277 (.A1(I355), .A2(I2379), .ZN(W277));
	NANDX1 U278 (.A1(I32), .A2(I65), .ZN(W278));
	NOR2X1 U281 (.A1(I3946), .A2(I410), .ZN(O129));
	INVX1 U282 (.I(I849), .ZN(O65));
	NANDX1 U284 (.A1(O381), .A2(I3958), .ZN(W284));
	NANDX1 U285 (.A1(I2784), .A2(I1961), .ZN(W285));
	NOR2X1 U289 (.A1(I1234), .A2(I1387), .ZN(W289));
	NANDX1 U297 (.A1(I1966), .A2(I50), .ZN(W297));
	NOR2X1 U303 (.A1(I2726), .A2(I4320), .ZN(W303));
	NANDX1 U304 (.A1(I953), .A2(I273), .ZN(W304));
	NOR2X1 U305 (.A1(O330), .A2(I2448), .ZN(W305));
	NANDX1 U306 (.A1(I4257), .A2(I1171), .ZN(W306));
	NOR2X1 U307 (.A1(I3655), .A2(I3116), .ZN(O179));
	INVX1 U311 (.I(I2654), .ZN(W311));
	NOR2X1 U318 (.A1(I3041), .A2(O65), .ZN(W318));
	NOR2X1 U319 (.A1(I981), .A2(I36), .ZN(W319));
	INVX1 U322 (.I(I2464), .ZN(W322));
	NANDX1 U323 (.A1(I1976), .A2(I2422), .ZN(W323));
	NOR2X1 U324 (.A1(W207), .A2(I2790), .ZN(W324));
	INVX1 U325 (.I(I453), .ZN(W325));
	INVX1 U327 (.I(I680), .ZN(W327));
	NANDX1 U330 (.A1(I940), .A2(I2598), .ZN(W330));
	NANDX1 U335 (.A1(I4338), .A2(I3523), .ZN(O173));
	INVX1 U336 (.I(I690), .ZN(W336));
	INVX1 U341 (.I(I4619), .ZN(W341));
	INVX1 U344 (.I(I2588), .ZN(W344));
	NOR2X1 U345 (.A1(W289), .A2(I1798), .ZN(W345));
	INVX1 U347 (.I(I3888), .ZN(W347));
	NOR2X1 U352 (.A1(I4990), .A2(I3302), .ZN(W352));
	INVX1 U355 (.I(I1489), .ZN(W355));
	INVX1 U357 (.I(I2034), .ZN(W357));
	NOR2X1 U358 (.A1(I216), .A2(I833), .ZN(W358));
	NOR2X1 U360 (.A1(I4367), .A2(I4662), .ZN(W360));
	NANDX1 U369 (.A1(I1481), .A2(I292), .ZN(O81));
	INVX1 U370 (.I(I107), .ZN(W370));
	NOR2X1 U374 (.A1(I3014), .A2(I4341), .ZN(W374));
	NANDX1 U378 (.A1(I404), .A2(I3516), .ZN(W378));
	INVX1 U382 (.I(I831), .ZN(W382));
	NANDX1 U388 (.A1(I1307), .A2(I2071), .ZN(W388));
	NOR2X1 U391 (.A1(I2919), .A2(I2939), .ZN(W391));
	INVX1 U394 (.I(I537), .ZN(W394));
	NOR2X1 U398 (.A1(I4268), .A2(I2957), .ZN(W398));
	INVX1 U400 (.I(I4039), .ZN(W400));
	INVX1 U404 (.I(I3312), .ZN(W404));
	NOR2X1 U405 (.A1(I1893), .A2(I3181), .ZN(W405));
	NOR2X1 U408 (.A1(I3206), .A2(I4174), .ZN(W408));
	NOR2X1 U409 (.A1(I1809), .A2(I1386), .ZN(W409));
	INVX1 U411 (.I(W311), .ZN(W411));
	NANDX1 U413 (.A1(I4325), .A2(I3213), .ZN(O428));
	NOR2X1 U414 (.A1(I4653), .A2(I3033), .ZN(W414));
	NOR2X1 U418 (.A1(I2132), .A2(I2191), .ZN(W418));
	NANDX1 U419 (.A1(I674), .A2(I3658), .ZN(W419));
	NANDX1 U423 (.A1(I3999), .A2(I2144), .ZN(W423));
	NOR2X1 U424 (.A1(I2453), .A2(W112), .ZN(W424));
	INVX1 U426 (.I(I3722), .ZN(W426));
	INVX1 U428 (.I(W50), .ZN(W428));
	NOR2X1 U430 (.A1(W388), .A2(O129), .ZN(W430));
	NOR2X1 U432 (.A1(W215), .A2(I2863), .ZN(W432));
	INVX1 U433 (.I(I4939), .ZN(W433));
	NOR2X1 U434 (.A1(I2466), .A2(I2342), .ZN(O197));
	NANDX1 U437 (.A1(I578), .A2(W5), .ZN(W437));
	INVX1 U440 (.I(W360), .ZN(W440));
	NOR2X1 U441 (.A1(I2513), .A2(I674), .ZN(W441));
	NOR2X1 U442 (.A1(I1130), .A2(I4908), .ZN(W442));
	NANDX1 U445 (.A1(I2612), .A2(I1221), .ZN(W445));
	INVX1 U446 (.I(I1176), .ZN(W446));
	NANDX1 U447 (.A1(W58), .A2(I3118), .ZN(W447));
	NOR2X1 U449 (.A1(W96), .A2(I638), .ZN(W449));
	NOR2X1 U450 (.A1(I3590), .A2(I2687), .ZN(W450));
	INVX1 U451 (.I(I4103), .ZN(W451));
	NANDX1 U453 (.A1(I2775), .A2(I996), .ZN(W453));
	INVX1 U456 (.I(I2268), .ZN(W456));
	INVX1 U458 (.I(W140), .ZN(W458));
	NANDX1 U459 (.A1(I3789), .A2(I2463), .ZN(W459));
	NANDX1 U463 (.A1(I1519), .A2(I3594), .ZN(W463));
	NANDX1 U466 (.A1(I4393), .A2(I33), .ZN(W466));
	INVX1 U468 (.I(I681), .ZN(W468));
	NOR2X1 U470 (.A1(I3245), .A2(I766), .ZN(W470));
	NOR2X1 U471 (.A1(I261), .A2(I3229), .ZN(W471));
	NANDX1 U476 (.A1(I1549), .A2(I4537), .ZN(W476));
	NOR2X1 U479 (.A1(I1346), .A2(I3777), .ZN(W479));
	NANDX1 U481 (.A1(I2319), .A2(W199), .ZN(W481));
	NANDX1 U486 (.A1(W453), .A2(I4017), .ZN(W486));
	NOR2X1 U487 (.A1(I3506), .A2(I1351), .ZN(W487));
	INVX1 U488 (.I(I4063), .ZN(W488));
	NOR2X1 U493 (.A1(I1534), .A2(I1756), .ZN(W493));
	INVX1 U497 (.I(I4313), .ZN(W497));
	NANDX1 U498 (.A1(I1772), .A2(I1653), .ZN(W498));
	INVX1 U499 (.I(I1249), .ZN(W499));
	INVX1 U504 (.I(I1976), .ZN(W504));
	INVX1 U507 (.I(W400), .ZN(O244));
	INVX1 U510 (.I(W180), .ZN(W510));
	INVX1 U513 (.I(W437), .ZN(W513));
	NOR2X1 U515 (.A1(I4217), .A2(I4671), .ZN(W515));
	INVX1 U516 (.I(I648), .ZN(W516));
	INVX1 U517 (.I(W264), .ZN(W517));
	NOR2X1 U519 (.A1(I4415), .A2(I1609), .ZN(W519));
	NANDX1 U526 (.A1(I187), .A2(I3548), .ZN(W526));
	INVX1 U528 (.I(I4436), .ZN(W528));
	INVX1 U529 (.I(I2237), .ZN(W529));
	NANDX1 U530 (.A1(I2304), .A2(I746), .ZN(O334));
	INVX1 U531 (.I(I4008), .ZN(W531));
	INVX1 U533 (.I(I1922), .ZN(W533));
	NOR2X1 U534 (.A1(I1162), .A2(I3081), .ZN(W534));
	NOR2X1 U536 (.A1(I823), .A2(I1146), .ZN(W536));
	NANDX1 U537 (.A1(W318), .A2(I549), .ZN(W537));
	NANDX1 U541 (.A1(I669), .A2(I3301), .ZN(W541));
	NOR2X1 U544 (.A1(W120), .A2(I1082), .ZN(O378));
	NANDX1 U547 (.A1(I2835), .A2(O65), .ZN(W547));
	NANDX1 U548 (.A1(I2229), .A2(I3305), .ZN(W548));
	NOR2X1 U556 (.A1(I4534), .A2(I777), .ZN(W556));
	INVX1 U564 (.I(W212), .ZN(W564));
	NOR2X1 U565 (.A1(I4534), .A2(I3354), .ZN(W565));
	INVX1 U568 (.I(W72), .ZN(W568));
	NANDX1 U569 (.A1(I1838), .A2(I1947), .ZN(O15));
	NANDX1 U571 (.A1(I4710), .A2(I2001), .ZN(W571));
	NOR2X1 U572 (.A1(I1473), .A2(W63), .ZN(O211));
	NOR2X1 U575 (.A1(W468), .A2(I878), .ZN(W575));
	INVX1 U577 (.I(I4351), .ZN(W577));
	NANDX1 U581 (.A1(I1670), .A2(I3606), .ZN(W581));
	INVX1 U582 (.I(I4925), .ZN(W582));
	NANDX1 U585 (.A1(I481), .A2(I2359), .ZN(W585));
	NANDX1 U589 (.A1(I2836), .A2(I4043), .ZN(W589));
	INVX1 U593 (.I(W515), .ZN(W593));
	INVX1 U595 (.I(W341), .ZN(W595));
	INVX1 U596 (.I(I3286), .ZN(W596));
	NOR2X1 U599 (.A1(I713), .A2(I2637), .ZN(W599));
	NANDX1 U600 (.A1(W63), .A2(I142), .ZN(W600));
	INVX1 U603 (.I(I3293), .ZN(W603));
	NANDX1 U604 (.A1(I4952), .A2(I72), .ZN(W604));
	NANDX1 U606 (.A1(W91), .A2(I565), .ZN(W606));
	NOR2X1 U607 (.A1(W327), .A2(I4795), .ZN(W607));
	NANDX1 U614 (.A1(W102), .A2(I4107), .ZN(W614));
	INVX1 U616 (.I(I2413), .ZN(O336));
	NOR2X1 U617 (.A1(I3070), .A2(I2310), .ZN(W617));
	NANDX1 U619 (.A1(I1303), .A2(I134), .ZN(W619));
	INVX1 U621 (.I(I4119), .ZN(W621));
	NANDX1 U624 (.A1(I3610), .A2(I3416), .ZN(W624));
	NANDX1 U625 (.A1(W437), .A2(I4850), .ZN(W625));
	NOR2X1 U626 (.A1(I4131), .A2(I2562), .ZN(W626));
	NOR2X1 U630 (.A1(I4127), .A2(I461), .ZN(W630));
	NANDX1 U631 (.A1(I3266), .A2(I1688), .ZN(W631));
	INVX1 U632 (.I(I1040), .ZN(O172));
	NANDX1 U633 (.A1(I2397), .A2(I1150), .ZN(W633));
	NOR2X1 U634 (.A1(I3367), .A2(I4129), .ZN(W634));
	INVX1 U635 (.I(I2531), .ZN(W635));
	NANDX1 U637 (.A1(I4409), .A2(I4269), .ZN(W637));
	NOR2X1 U638 (.A1(I2124), .A2(I2350), .ZN(W638));
	INVX1 U639 (.I(I3157), .ZN(W639));
	INVX1 U640 (.I(I849), .ZN(W640));
	NANDX1 U642 (.A1(I2539), .A2(W53), .ZN(W642));
	NOR2X1 U645 (.A1(W330), .A2(I2975), .ZN(O467));
	NOR2X1 U646 (.A1(W278), .A2(I3843), .ZN(W646));
	INVX1 U649 (.I(I4003), .ZN(W649));
	NANDX1 U652 (.A1(W577), .A2(I2583), .ZN(W652));
	NANDX1 U660 (.A1(I1690), .A2(I3109), .ZN(W660));
	INVX1 U661 (.I(I891), .ZN(W661));
	NOR2X1 U664 (.A1(I3208), .A2(W355), .ZN(W664));
	NANDX1 U665 (.A1(W69), .A2(I1931), .ZN(W665));
	NANDX1 U667 (.A1(O296), .A2(I3529), .ZN(W667));
	NOR2X1 U669 (.A1(I3301), .A2(I3309), .ZN(O411));
	INVX1 U671 (.I(I1936), .ZN(W671));
	NANDX1 U672 (.A1(I3245), .A2(I1678), .ZN(O191));
	NANDX1 U674 (.A1(I1929), .A2(I262), .ZN(W674));
	NANDX1 U676 (.A1(I4132), .A2(I4993), .ZN(W676));
	INVX1 U677 (.I(I1462), .ZN(O180));
	INVX1 U683 (.I(I1712), .ZN(W683));
	NANDX1 U686 (.A1(I548), .A2(W138), .ZN(W686));
	NANDX1 U691 (.A1(W589), .A2(I1805), .ZN(W691));
	NANDX1 U693 (.A1(W74), .A2(I3234), .ZN(W693));
	NOR2X1 U696 (.A1(I1387), .A2(I377), .ZN(O346));
	INVX1 U697 (.I(W90), .ZN(W697));
	NANDX1 U702 (.A1(I1128), .A2(I2361), .ZN(W702));
	NANDX1 U707 (.A1(I2019), .A2(I4545), .ZN(W707));
	NOR2X1 U710 (.A1(I1834), .A2(I3187), .ZN(O433));
	NANDX1 U711 (.A1(I1097), .A2(I2187), .ZN(W711));
	INVX1 U712 (.I(I845), .ZN(W712));
	INVX1 U713 (.I(I337), .ZN(W713));
	INVX1 U716 (.I(I1150), .ZN(W716));
	INVX1 U720 (.I(W153), .ZN(W720));
	INVX1 U721 (.I(I2349), .ZN(O459));
	NOR2X1 U722 (.A1(I1639), .A2(W303), .ZN(O359));
	INVX1 U723 (.I(I3896), .ZN(O288));
	NOR2X1 U728 (.A1(I4090), .A2(I3885), .ZN(W728));
	INVX1 U729 (.I(I3621), .ZN(W729));
	NANDX1 U731 (.A1(I1401), .A2(I3519), .ZN(W731));
	NANDX1 U735 (.A1(I1174), .A2(I2566), .ZN(W735));
	INVX1 U745 (.I(I1808), .ZN(W745));
	NANDX1 U746 (.A1(I213), .A2(I2743), .ZN(O377));
	NOR2X1 U747 (.A1(I41), .A2(W153), .ZN(W747));
	NANDX1 U748 (.A1(I3007), .A2(I2313), .ZN(W748));
	NOR2X1 U750 (.A1(W166), .A2(I650), .ZN(W750));
	INVX1 U751 (.I(W638), .ZN(O385));
	NOR2X1 U756 (.A1(I3707), .A2(I880), .ZN(W756));
	NOR2X1 U757 (.A1(I878), .A2(I4081), .ZN(W757));
	INVX1 U759 (.I(I1410), .ZN(W759));
	NOR2X1 U760 (.A1(I2944), .A2(I2644), .ZN(W760));
	INVX1 U764 (.I(I3019), .ZN(W764));
	NOR2X1 U766 (.A1(I1291), .A2(I3401), .ZN(W766));
	INVX1 U770 (.I(I1805), .ZN(O282));
	NOR2X1 U771 (.A1(I3875), .A2(I4877), .ZN(W771));
	NANDX1 U775 (.A1(I1605), .A2(I1314), .ZN(W775));
	INVX1 U776 (.I(I717), .ZN(W776));
	INVX1 U781 (.I(I731), .ZN(O395));
	NANDX1 U782 (.A1(I639), .A2(I960), .ZN(W782));
	NOR2X1 U783 (.A1(O378), .A2(I2561), .ZN(W783));
	NANDX1 U784 (.A1(I2404), .A2(I2513), .ZN(W784));
	INVX1 U785 (.I(I393), .ZN(W785));
	INVX1 U786 (.I(I4906), .ZN(W786));
	INVX1 U787 (.I(I3095), .ZN(W787));
	NANDX1 U788 (.A1(W404), .A2(I4083), .ZN(W788));
	NANDX1 U791 (.A1(I4784), .A2(I4480), .ZN(W791));
	NANDX1 U792 (.A1(I3787), .A2(I3732), .ZN(W792));
	INVX1 U796 (.I(W526), .ZN(W796));
	INVX1 U797 (.I(I846), .ZN(W797));
	NANDX1 U800 (.A1(W440), .A2(I17), .ZN(W800));
	NANDX1 U802 (.A1(I1589), .A2(I3540), .ZN(W802));
	NANDX1 U803 (.A1(W449), .A2(W720), .ZN(W803));
	NANDX1 U805 (.A1(W352), .A2(I1009), .ZN(W805));
	NANDX1 U807 (.A1(I1893), .A2(I482), .ZN(W807));
	NANDX1 U808 (.A1(W325), .A2(I252), .ZN(O311));
	NOR2X1 U811 (.A1(I1000), .A2(W246), .ZN(W811));
	INVX1 U817 (.I(I3232), .ZN(O253));
	NANDX1 U819 (.A1(I3355), .A2(W374), .ZN(O219));
	NANDX1 U826 (.A1(I1306), .A2(I1547), .ZN(W826));
	INVX1 U831 (.I(W306), .ZN(W831));
	INVX1 U832 (.I(I903), .ZN(O47));
	INVX1 U833 (.I(I3901), .ZN(W833));
	NANDX1 U837 (.A1(O288), .A2(I4807), .ZN(W837));
	NANDX1 U838 (.A1(W411), .A2(I2673), .ZN(W838));
	NANDX1 U840 (.A1(W716), .A2(I2880), .ZN(W840));
	INVX1 U841 (.I(I1438), .ZN(W841));
	NOR2X1 U842 (.A1(I1266), .A2(I3594), .ZN(W842));
	INVX1 U848 (.I(I937), .ZN(W848));
	NANDX1 U854 (.A1(I3567), .A2(I2498), .ZN(W854));
	NANDX1 U856 (.A1(I1089), .A2(W614), .ZN(W856));
	NOR2X1 U860 (.A1(W488), .A2(I598), .ZN(W860));
	NOR2X1 U864 (.A1(W671), .A2(W831), .ZN(W864));
	NOR2X1 U869 (.A1(I618), .A2(I3167), .ZN(W869));
	NOR2X1 U873 (.A1(I2420), .A2(I3160), .ZN(W873));
	NANDX1 U878 (.A1(I2360), .A2(I1846), .ZN(W878));
	INVX1 U879 (.I(I548), .ZN(W879));
	NOR2X1 U881 (.A1(I4791), .A2(I928), .ZN(W881));
	INVX1 U882 (.I(W660), .ZN(W882));
	NOR2X1 U884 (.A1(W881), .A2(I4291), .ZN(W884));
	NOR2X1 U885 (.A1(W39), .A2(I4288), .ZN(W885));
	INVX1 U888 (.I(I1186), .ZN(W888));
	INVX1 U890 (.I(I232), .ZN(W890));
	NOR2X1 U896 (.A1(O173), .A2(W11), .ZN(W896));
	NOR2X1 U897 (.A1(I3629), .A2(I4815), .ZN(O181));
	NANDX1 U898 (.A1(I1455), .A2(I218), .ZN(W898));
	NANDX1 U899 (.A1(I2413), .A2(I1094), .ZN(W899));
	INVX1 U900 (.I(I1043), .ZN(O406));
	INVX1 U901 (.I(W513), .ZN(W901));
	INVX1 U902 (.I(W805), .ZN(W902));
	INVX1 U904 (.I(I4211), .ZN(W904));
	NOR2X1 U905 (.A1(I3941), .A2(I1855), .ZN(O152));
	INVX1 U908 (.I(I4597), .ZN(W908));
	INVX1 U909 (.I(I850), .ZN(W909));
	INVX1 U913 (.I(I644), .ZN(W913));
	INVX1 U914 (.I(I3848), .ZN(W914));
	NANDX1 U915 (.A1(W493), .A2(I319), .ZN(W915));
	INVX1 U918 (.I(W712), .ZN(W918));
	INVX1 U924 (.I(I1579), .ZN(W924));
	NOR2X1 U926 (.A1(I2614), .A2(I453), .ZN(W926));
	NANDX1 U929 (.A1(I506), .A2(I4170), .ZN(W929));
	NANDX1 U932 (.A1(W479), .A2(W126), .ZN(W932));
	NANDX1 U935 (.A1(W785), .A2(I123), .ZN(W935));
	INVX1 U936 (.I(I674), .ZN(O283));
	NANDX1 U942 (.A1(I431), .A2(I4829), .ZN(W942));
	INVX1 U943 (.I(W826), .ZN(O458));
	NOR2X1 U944 (.A1(I3565), .A2(I2953), .ZN(W944));
	NOR2X1 U948 (.A1(I3233), .A2(I1891), .ZN(O162));
	NOR2X1 U952 (.A1(I1086), .A2(W792), .ZN(W952));
	NANDX1 U954 (.A1(I602), .A2(I818), .ZN(W954));
	NANDX1 U957 (.A1(I3984), .A2(I1354), .ZN(W957));
	NOR2X1 U959 (.A1(I2809), .A2(I904), .ZN(W959));
	NOR2X1 U960 (.A1(I3390), .A2(I4337), .ZN(W960));
	NOR2X1 U961 (.A1(I4642), .A2(I63), .ZN(O183));
	NANDX1 U964 (.A1(I4253), .A2(I1101), .ZN(W964));
	INVX1 U972 (.I(W683), .ZN(W972));
	NANDX1 U973 (.A1(I2786), .A2(I474), .ZN(W973));
	INVX1 U976 (.I(I3021), .ZN(W976));
	NANDX1 U977 (.A1(O172), .A2(I895), .ZN(W977));
	NANDX1 U980 (.A1(I3738), .A2(I3293), .ZN(W980));
	INVX1 U982 (.I(I630), .ZN(W982));
	NOR2X1 U983 (.A1(I2717), .A2(I2189), .ZN(W983));
	NOR2X1 U984 (.A1(W144), .A2(W631), .ZN(W984));
	INVX1 U985 (.I(W944), .ZN(W985));
	NOR2X1 U987 (.A1(I2639), .A2(W756), .ZN(W987));
	NANDX1 U988 (.A1(I4376), .A2(W217), .ZN(W988));
	NANDX1 U991 (.A1(I3384), .A2(I1403), .ZN(W991));
	NOR2X1 U992 (.A1(O136), .A2(I700), .ZN(W992));
	INVX1 U993 (.I(I2504), .ZN(O79));
	NOR2X1 U1000 (.A1(W265), .A2(I370), .ZN(O420));
	NOR2X1 U1002 (.A1(I4826), .A2(W201), .ZN(W1002));
	NOR2X1 U1003 (.A1(I2622), .A2(I2667), .ZN(O241));
	NANDX1 U1004 (.A1(I66), .A2(I4961), .ZN(W1004));
	NOR2X1 U1012 (.A1(I1226), .A2(I3738), .ZN(W1012));
	INVX1 U1014 (.I(W344), .ZN(W1014));
	NANDX1 U1016 (.A1(W382), .A2(O296), .ZN(W1016));
	INVX1 U1018 (.I(I3991), .ZN(O441));
	NANDX1 U1019 (.A1(W757), .A2(I3269), .ZN(W1019));
	NOR2X1 U1026 (.A1(I2069), .A2(W848), .ZN(W1026));
	NOR2X1 U1027 (.A1(I1031), .A2(I2192), .ZN(W1027));
	INVX1 U1028 (.I(I1813), .ZN(W1028));
	NANDX1 U1033 (.A1(I2540), .A2(I950), .ZN(W1033));
	NOR2X1 U1036 (.A1(I1724), .A2(W621), .ZN(W1036));
	NANDX1 U1037 (.A1(I241), .A2(W957), .ZN(W1037));
	NANDX1 U1038 (.A1(W841), .A2(W305), .ZN(W1038));
	NOR2X1 U1039 (.A1(I3153), .A2(I2877), .ZN(W1039));
	NOR2X1 U1040 (.A1(I726), .A2(W504), .ZN(W1040));
	NANDX1 U1043 (.A1(W107), .A2(I2295), .ZN(O91));
	INVX1 U1044 (.I(I2682), .ZN(W1044));
	INVX1 U1045 (.I(W414), .ZN(W1045));
	INVX1 U1048 (.I(I1189), .ZN(W1048));
	INVX1 U1050 (.I(I162), .ZN(W1050));
	NANDX1 U1059 (.A1(I2294), .A2(W1004), .ZN(W1059));
	NANDX1 U1061 (.A1(I2406), .A2(W1038), .ZN(W1061));
	INVX1 U1064 (.I(I4414), .ZN(W1064));
	NANDX1 U1065 (.A1(W879), .A2(W8), .ZN(W1065));
	INVX1 U1066 (.I(W571), .ZN(W1066));
	NOR2X1 U1067 (.A1(I3039), .A2(I2495), .ZN(W1067));
	INVX1 U1069 (.I(I2061), .ZN(W1069));
	INVX1 U1071 (.I(I375), .ZN(O68));
	NANDX1 U1079 (.A1(W599), .A2(W926), .ZN(W1079));
	NANDX1 U1085 (.A1(I32), .A2(W456), .ZN(W1085));
	NANDX1 U1091 (.A1(I2349), .A2(O482), .ZN(W1091));
	NANDX1 U1092 (.A1(I2303), .A2(I2277), .ZN(W1092));
	NANDX1 U1095 (.A1(I310), .A2(W510), .ZN(W1095));
	NOR2X1 U1096 (.A1(W884), .A2(I3959), .ZN(W1096));
	INVX1 U1097 (.I(W423), .ZN(W1097));
	NOR2X1 U1108 (.A1(I1266), .A2(I2018), .ZN(W1108));
	NANDX1 U1113 (.A1(I1314), .A2(I36), .ZN(W1113));
	INVX1 U1117 (.I(I444), .ZN(W1117));
	NANDX1 U1118 (.A1(W918), .A2(W954), .ZN(W1118));
	NOR2X1 U1120 (.A1(I303), .A2(I4848), .ZN(W1120));
	INVX1 U1125 (.I(W833), .ZN(O147));
	NOR2X1 U1126 (.A1(W756), .A2(W537), .ZN(W1126));
	NOR2X1 U1132 (.A1(I3266), .A2(I3633), .ZN(O478));
	NANDX1 U1133 (.A1(I532), .A2(W107), .ZN(W1133));
	INVX1 U1135 (.I(I787), .ZN(O196));
	NANDX1 U1138 (.A1(W759), .A2(I3195), .ZN(W1138));
	NANDX1 U1139 (.A1(W319), .A2(I4339), .ZN(W1139));
	NOR2X1 U1140 (.A1(W1139), .A2(I3363), .ZN(W1140));
	NANDX1 U1145 (.A1(W198), .A2(I2446), .ZN(W1145));
	INVX1 U1147 (.I(W1133), .ZN(O165));
	NOR2X1 U1149 (.A1(W113), .A2(I4103), .ZN(O146));
	INVX1 U1151 (.I(W984), .ZN(O369));
	NANDX1 U1153 (.A1(I2238), .A2(I1575), .ZN(W1153));
	NANDX1 U1154 (.A1(I749), .A2(I833), .ZN(W1154));
	NANDX1 U1158 (.A1(I970), .A2(I3709), .ZN(W1158));
	INVX1 U1160 (.I(I3507), .ZN(W1160));
	INVX1 U1168 (.I(W1002), .ZN(W1168));
	NANDX1 U1172 (.A1(W155), .A2(I2968), .ZN(W1172));
	INVX1 U1178 (.I(W285), .ZN(W1178));
	NANDX1 U1179 (.A1(I1443), .A2(I398), .ZN(W1179));
	NANDX1 U1182 (.A1(I3497), .A2(I1533), .ZN(W1182));
	INVX1 U1185 (.I(I4713), .ZN(W1185));
	INVX1 U1186 (.I(I1497), .ZN(W1186));
	NANDX1 U1188 (.A1(I4530), .A2(W1079), .ZN(W1188));
	NOR2X1 U1189 (.A1(O482), .A2(W336), .ZN(W1189));
	NOR2X1 U1190 (.A1(I3013), .A2(W360), .ZN(W1190));
	NANDX1 U1192 (.A1(I4654), .A2(I499), .ZN(W1192));
	NOR2X1 U1194 (.A1(I4660), .A2(I3519), .ZN(W1194));
	NANDX1 U1195 (.A1(I174), .A2(I2000), .ZN(O422));
	INVX1 U1196 (.I(W114), .ZN(O209));
	NANDX1 U1201 (.A1(I3092), .A2(I1051), .ZN(W1201));
	NOR2X1 U1205 (.A1(I4803), .A2(I2309), .ZN(W1205));
	NANDX1 U1206 (.A1(W533), .A2(I2544), .ZN(O61));
	INVX1 U1211 (.I(W193), .ZN(W1211));
	INVX1 U1214 (.I(I4475), .ZN(W1214));
	NANDX1 U1216 (.A1(I3928), .A2(I3720), .ZN(W1216));
	INVX1 U1218 (.I(W987), .ZN(W1218));
	INVX1 U1219 (.I(W304), .ZN(W1219));
	NANDX1 U1225 (.A1(I3162), .A2(I956), .ZN(W1225));
	NOR2X1 U1231 (.A1(W581), .A2(I299), .ZN(W1231));
	NOR2X1 U1233 (.A1(I1565), .A2(I3334), .ZN(W1233));
	INVX1 U1234 (.I(I974), .ZN(W1234));
	INVX1 U1237 (.I(W17), .ZN(W1237));
	NANDX1 U1241 (.A1(I4112), .A2(W635), .ZN(W1241));
	INVX1 U1242 (.I(I3289), .ZN(W1242));
	INVX1 U1247 (.I(I1972), .ZN(W1247));
	NOR2X1 U1251 (.A1(I1944), .A2(I3727), .ZN(W1251));
	NOR2X1 U1253 (.A1(W106), .A2(I1137), .ZN(W1253));
	NOR2X1 U1263 (.A1(I260), .A2(I3623), .ZN(O333));
	INVX1 U1264 (.I(I1294), .ZN(O74));
	NANDX1 U1266 (.A1(I719), .A2(W776), .ZN(O265));
	INVX1 U1271 (.I(I3826), .ZN(O246));
	INVX1 U1272 (.I(W565), .ZN(W1272));
	NOR2X1 U1273 (.A1(I3528), .A2(W85), .ZN(W1273));
	NANDX1 U1274 (.A1(W973), .A2(W1012), .ZN(W1274));
	NOR2X1 U1275 (.A1(I3970), .A2(I3965), .ZN(W1275));
	NANDX1 U1284 (.A1(I1123), .A2(W890), .ZN(W1284));
	INVX1 U1285 (.I(I3890), .ZN(W1285));
	NOR2X1 U1286 (.A1(I2694), .A2(I1157), .ZN(O161));
	NOR2X1 U1289 (.A1(I2355), .A2(W391), .ZN(W1289));
	NANDX1 U1291 (.A1(W98), .A2(W1218), .ZN(W1291));
	INVX1 U1292 (.I(W129), .ZN(W1292));
	NOR2X1 U1293 (.A1(W661), .A2(I3381), .ZN(W1293));
	INVX1 U1297 (.I(I1783), .ZN(W1297));
	INVX1 U1300 (.I(I3314), .ZN(O319));
	NOR2X1 U1301 (.A1(I3003), .A2(I53), .ZN(W1301));
	INVX1 U1304 (.I(I2245), .ZN(W1304));
	INVX1 U1305 (.I(W547), .ZN(O276));
	NANDX1 U1311 (.A1(I385), .A2(I228), .ZN(W1311));
	NOR2X1 U1319 (.A1(I3974), .A2(I2568), .ZN(W1319));
	NANDX1 U1320 (.A1(I2874), .A2(W73), .ZN(W1320));
	NANDX1 U1322 (.A1(O420), .A2(I1272), .ZN(W1322));
	INVX1 U1324 (.I(W913), .ZN(W1324));
	INVX1 U1326 (.I(W69), .ZN(W1326));
	NOR2X1 U1328 (.A1(I1134), .A2(W697), .ZN(W1328));
	INVX1 U1329 (.I(I2357), .ZN(W1329));
	INVX1 U1331 (.I(I1668), .ZN(O141));
	NANDX1 U1334 (.A1(W1241), .A2(I652), .ZN(W1334));
	NANDX1 U1339 (.A1(I2077), .A2(W838), .ZN(W1339));
	NANDX1 U1341 (.A1(I3685), .A2(I1879), .ZN(W1341));
	INVX1 U1344 (.I(W782), .ZN(W1344));
	NOR2X1 U1345 (.A1(W924), .A2(W976), .ZN(W1345));
	NOR2X1 U1347 (.A1(W166), .A2(I2132), .ZN(O394));
	NOR2X1 U1350 (.A1(I87), .A2(I4177), .ZN(O460));
	NOR2X1 U1351 (.A1(I353), .A2(I3050), .ZN(W1351));
	NOR2X1 U1353 (.A1(I1202), .A2(I4785), .ZN(W1353));
	NANDX1 U1357 (.A1(I1308), .A2(W94), .ZN(W1357));
	INVX1 U1363 (.I(I1497), .ZN(W1363));
	NANDX1 U1370 (.A1(I3752), .A2(I4474), .ZN(W1370));
	NANDX1 U1372 (.A1(I3246), .A2(I2412), .ZN(W1372));
	NANDX1 U1373 (.A1(I4750), .A2(W642), .ZN(W1373));
	NANDX1 U1374 (.A1(I2885), .A2(I931), .ZN(W1374));
	NANDX1 U1377 (.A1(W1231), .A2(W942), .ZN(W1377));
	NOR2X1 U1380 (.A1(I2649), .A2(I4205), .ZN(W1380));
	NOR2X1 U1381 (.A1(W667), .A2(I4434), .ZN(W1381));
	INVX1 U1382 (.I(W357), .ZN(W1382));
	NOR2X1 U1386 (.A1(W1201), .A2(W161), .ZN(W1386));
	NOR2X1 U1387 (.A1(I4090), .A2(W599), .ZN(W1387));
	INVX1 U1388 (.I(I623), .ZN(W1388));
	NANDX1 U1389 (.A1(I347), .A2(I341), .ZN(W1389));
	NOR2X1 U1392 (.A1(I3067), .A2(W1334), .ZN(W1392));
	NANDX1 U1394 (.A1(W529), .A2(I934), .ZN(O335));
	NANDX1 U1396 (.A1(I2264), .A2(I3396), .ZN(W1396));
	NOR2X1 U1399 (.A1(I4488), .A2(I527), .ZN(W1399));
	INVX1 U1400 (.I(I4608), .ZN(W1400));
	NANDX1 U1401 (.A1(W1117), .A2(I3351), .ZN(W1401));
	NANDX1 U1405 (.A1(W646), .A2(I382), .ZN(W1405));
	NANDX1 U1408 (.A1(I4336), .A2(I4689), .ZN(W1408));
	NANDX1 U1410 (.A1(I1098), .A2(W497), .ZN(W1410));
	NOR2X1 U1411 (.A1(I584), .A2(I2533), .ZN(W1411));
	NOR2X1 U1415 (.A1(W152), .A2(I2687), .ZN(W1415));
	INVX1 U1416 (.I(I866), .ZN(W1416));
	NANDX1 U1417 (.A1(I1595), .A2(I2803), .ZN(W1417));
	INVX1 U1420 (.I(I349), .ZN(W1420));
	INVX1 U1425 (.I(I3032), .ZN(W1425));
	NANDX1 U1426 (.A1(I4152), .A2(W114), .ZN(O259));
	INVX1 U1430 (.I(I147), .ZN(W1430));
	INVX1 U1433 (.I(I4133), .ZN(W1433));
	NANDX1 U1434 (.A1(I3390), .A2(I1008), .ZN(W1434));
	INVX1 U1439 (.I(W1065), .ZN(W1439));
	NOR2X1 U1454 (.A1(W1411), .A2(W985), .ZN(W1454));
	NOR2X1 U1455 (.A1(I3381), .A2(W1326), .ZN(O114));
	INVX1 U1458 (.I(I4584), .ZN(W1458));
	NOR2X1 U1462 (.A1(I2884), .A2(I2904), .ZN(W1462));
	NANDX1 U1469 (.A1(I3507), .A2(I2098), .ZN(W1469));
	NANDX1 U1470 (.A1(W1059), .A2(I3252), .ZN(W1470));
	INVX1 U1473 (.I(W1092), .ZN(W1473));
	NANDX1 U1474 (.A1(I407), .A2(W21), .ZN(W1474));
	INVX1 U1476 (.I(W1027), .ZN(W1476));
	NANDX1 U1477 (.A1(I819), .A2(W791), .ZN(W1477));
	NANDX1 U1482 (.A1(I2966), .A2(W1462), .ZN(W1482));
	INVX1 U1489 (.I(I4559), .ZN(W1489));
	NANDX1 U1490 (.A1(W497), .A2(W277), .ZN(W1490));
	NANDX1 U1493 (.A1(I4368), .A2(I2801), .ZN(O109));
	NANDX1 U1495 (.A1(I2630), .A2(I2752), .ZN(W1495));
	NOR2X1 U1496 (.A1(I3631), .A2(I2006), .ZN(W1496));
	NOR2X1 U1502 (.A1(I1353), .A2(I2302), .ZN(W1502));
	INVX1 U1503 (.I(O408), .ZN(W1503));
	INVX1 U1509 (.I(W633), .ZN(W1509));
	NOR2X1 U1517 (.A1(I2324), .A2(W40), .ZN(W1517));
	NOR2X1 U1519 (.A1(I3631), .A2(I4720), .ZN(W1519));
	INVX1 U1523 (.I(I1893), .ZN(W1523));
	NOR2X1 U1527 (.A1(W1085), .A2(W536), .ZN(W1527));
	NANDX1 U1528 (.A1(I1467), .A2(I1649), .ZN(W1528));
	NOR2X1 U1530 (.A1(I4852), .A2(I1366), .ZN(O227));
	NANDX1 U1536 (.A1(I3350), .A2(I3174), .ZN(W1536));
	NANDX1 U1537 (.A1(I3972), .A2(I3172), .ZN(W1537));
	INVX1 U1538 (.I(W531), .ZN(W1538));
	INVX1 U1539 (.I(I2822), .ZN(W1539));
	INVX1 U1540 (.I(W1399), .ZN(W1540));
	INVX1 U1541 (.I(O61), .ZN(W1541));
	NANDX1 U1547 (.A1(I4720), .A2(I1837), .ZN(O324));
	NANDX1 U1548 (.A1(I393), .A2(W510), .ZN(W1548));
	INVX1 U1558 (.I(I1754), .ZN(W1558));
	NANDX1 U1561 (.A1(W585), .A2(O72), .ZN(W1561));
	INVX1 U1562 (.I(W1061), .ZN(W1562));
	NOR2X1 U1564 (.A1(W1108), .A2(W1319), .ZN(W1564));
	NANDX1 U1566 (.A1(W1097), .A2(W1381), .ZN(W1566));
	NOR2X1 U1567 (.A1(W711), .A2(I3407), .ZN(W1567));
	NOR2X1 U1568 (.A1(W1251), .A2(I4836), .ZN(W1568));
	INVX1 U1571 (.I(I2523), .ZN(W1571));
	INVX1 U1573 (.I(I3724), .ZN(O185));
	NOR2X1 U1574 (.A1(I2922), .A2(W442), .ZN(W1574));
	NANDX1 U1581 (.A1(I3323), .A2(I437), .ZN(W1581));
	NOR2X1 U1585 (.A1(I4744), .A2(W964), .ZN(W1585));
	INVX1 U1586 (.I(I1466), .ZN(O215));
	INVX1 U1587 (.I(I3195), .ZN(O30));
	NANDX1 U1589 (.A1(I4282), .A2(I4280), .ZN(W1589));
	NOR2X1 U1592 (.A1(I642), .A2(W162), .ZN(W1592));
	NOR2X1 U1593 (.A1(I1244), .A2(I3341), .ZN(W1593));
	NANDX1 U1598 (.A1(I2589), .A2(W982), .ZN(W1598));
	NOR2X1 U1604 (.A1(I4686), .A2(W1489), .ZN(W1604));
	NANDX1 U1610 (.A1(I1244), .A2(I3683), .ZN(W1610));
	NANDX1 U1620 (.A1(I1031), .A2(I1562), .ZN(W1620));
	NANDX1 U1624 (.A1(I1734), .A2(I2402), .ZN(W1624));
	NANDX1 U1626 (.A1(I4902), .A2(I1500), .ZN(O21));
	INVX1 U1633 (.I(I1802), .ZN(W1633));
	INVX1 U1637 (.I(I2578), .ZN(W1637));
	INVX1 U1642 (.I(W1567), .ZN(W1642));
	NANDX1 U1652 (.A1(I256), .A2(W358), .ZN(O348));
	NOR2X1 U1655 (.A1(W1523), .A2(O215), .ZN(W1655));
	INVX1 U1656 (.I(W1192), .ZN(W1656));
	NOR2X1 U1657 (.A1(W973), .A2(I1369), .ZN(W1657));
	INVX1 U1659 (.I(I2724), .ZN(W1659));
	INVX1 U1661 (.I(I4247), .ZN(W1661));
	NOR2X1 U1668 (.A1(W667), .A2(I1214), .ZN(O192));
	NANDX1 U1672 (.A1(W1566), .A2(W433), .ZN(W1672));
	INVX1 U1673 (.I(W1118), .ZN(W1673));
	INVX1 U1679 (.I(I1814), .ZN(W1679));
	NOR2X1 U1680 (.A1(W1014), .A2(W634), .ZN(W1680));
	NANDX1 U1684 (.A1(I561), .A2(W1673), .ZN(O261));
	NANDX1 U1688 (.A1(I131), .A2(I3075), .ZN(W1688));
	INVX1 U1690 (.I(I3290), .ZN(W1690));
	NANDX1 U1691 (.A1(W398), .A2(I186), .ZN(W1691));
	NOR2X1 U1693 (.A1(I4714), .A2(I1721), .ZN(W1693));
	NANDX1 U1697 (.A1(I1576), .A2(I822), .ZN(W1697));
	NOR2X1 U1698 (.A1(W1377), .A2(W394), .ZN(W1698));
	NANDX1 U1704 (.A1(I4559), .A2(I1329), .ZN(O4));
	NOR2X1 U1714 (.A1(I3759), .A2(I3224), .ZN(W1714));
	NANDX1 U1718 (.A1(W860), .A2(I2306), .ZN(W1718));
	NANDX1 U1719 (.A1(W1108), .A2(W120), .ZN(W1719));
	NANDX1 U1720 (.A1(I51), .A2(I1218), .ZN(W1720));
	NOR2X1 U1721 (.A1(I1962), .A2(I1806), .ZN(W1721));
	NANDX1 U1725 (.A1(W47), .A2(W735), .ZN(W1725));
	INVX1 U1726 (.I(I1351), .ZN(W1726));
	INVX1 U1731 (.I(I3252), .ZN(O198));
	INVX1 U1732 (.I(W127), .ZN(W1732));
	NOR2X1 U1736 (.A1(W745), .A2(I4510), .ZN(W1736));
	INVX1 U1737 (.I(I4020), .ZN(W1737));
	NOR2X1 U1741 (.A1(W1726), .A2(W447), .ZN(W1741));
	NANDX1 U1742 (.A1(I1927), .A2(I2172), .ZN(W1742));
	NANDX1 U1743 (.A1(I3214), .A2(I2194), .ZN(O234));
	INVX1 U1744 (.I(I1641), .ZN(W1744));
	NANDX1 U1747 (.A1(I697), .A2(I2150), .ZN(W1747));
	INVX1 U1755 (.I(I3165), .ZN(O2));
	INVX1 U1761 (.I(W1016), .ZN(W1761));
	NANDX1 U1762 (.A1(I3360), .A2(I4618), .ZN(W1762));
	NOR2X1 U1763 (.A1(W516), .A2(W1231), .ZN(W1763));
	NANDX1 U1767 (.A1(I2916), .A2(W1069), .ZN(W1767));
	INVX1 U1769 (.I(W347), .ZN(W1769));
	NOR2X1 U1770 (.A1(I4304), .A2(W1598), .ZN(W1770));
	NOR2X1 U1772 (.A1(I4848), .A2(W1095), .ZN(W1772));
	NOR2X1 U1774 (.A1(I2664), .A2(W382), .ZN(W1774));
	NOR2X1 U1779 (.A1(W1691), .A2(I3035), .ZN(W1779));
	INVX1 U1781 (.I(I4010), .ZN(W1781));
	NOR2X1 U1785 (.A1(W1454), .A2(I255), .ZN(W1785));
	INVX1 U1795 (.I(W1140), .ZN(W1795));
	NANDX1 U1797 (.A1(W707), .A2(W1417), .ZN(W1797));
	NANDX1 U1799 (.A1(I2906), .A2(W1033), .ZN(W1799));
	NANDX1 U1801 (.A1(W652), .A2(I584), .ZN(W1801));
	INVX1 U1802 (.I(I741), .ZN(W1802));
	NOR2X1 U1806 (.A1(W517), .A2(I4794), .ZN(O187));
	NANDX1 U1811 (.A1(I3279), .A2(W954), .ZN(O491));
	NOR2X1 U1813 (.A1(W617), .A2(I1400), .ZN(W1813));
	INVX1 U1815 (.I(I4929), .ZN(W1815));
	NOR2X1 U1821 (.A1(W603), .A2(W1496), .ZN(W1821));
	INVX1 U1823 (.I(I2512), .ZN(W1823));
	NOR2X1 U1834 (.A1(I238), .A2(I1462), .ZN(W1834));
	INVX1 U1836 (.I(W1097), .ZN(O111));
	NOR2X1 U1837 (.A1(W873), .A2(I1914), .ZN(W1837));
	INVX1 U1838 (.I(O79), .ZN(O54));
	NOR2X1 U1839 (.A1(W497), .A2(W1113), .ZN(O73));
	NANDX1 U1841 (.A1(I2977), .A2(I3860), .ZN(O145));
	NOR2X1 U1844 (.A1(I4304), .A2(I4073), .ZN(W1844));
	INVX1 U1850 (.I(I3868), .ZN(W1850));
	INVX1 U1856 (.I(W1691), .ZN(O474));
	INVX1 U1861 (.I(W972), .ZN(O182));
	INVX1 U1863 (.I(I2249), .ZN(W1863));
	NANDX1 U1864 (.A1(W977), .A2(I795), .ZN(W1864));
	NANDX1 U1866 (.A1(W786), .A2(W797), .ZN(O424));
	NANDX1 U1867 (.A1(I2937), .A2(I139), .ZN(O132));
	INVX1 U1868 (.I(I723), .ZN(W1868));
	NOR2X1 U1869 (.A1(I3009), .A2(W1566), .ZN(O416));
	INVX1 U1874 (.I(W1785), .ZN(W1874));
	NANDX1 U1875 (.A1(I2148), .A2(I2465), .ZN(O475));
	NOR2X1 U1881 (.A1(W1864), .A2(I4775), .ZN(W1881));
	INVX1 U1886 (.I(I4464), .ZN(W1886));
	NOR2X1 U1890 (.A1(I4643), .A2(W74), .ZN(W1890));
	NANDX1 U1893 (.A1(I1369), .A2(I4698), .ZN(O176));
	NOR2X1 U1895 (.A1(I4924), .A2(W1581), .ZN(W1895));
	NANDX1 U1898 (.A1(I4036), .A2(I108), .ZN(O267));
	NOR2X1 U1906 (.A1(I4133), .A2(W479), .ZN(O299));
	NOR2X1 U1910 (.A1(W1291), .A2(W840), .ZN(W1910));
	INVX1 U1913 (.I(I2789), .ZN(W1913));
	NOR2X1 U1915 (.A1(I1480), .A2(W1844), .ZN(W1915));
	NOR2X1 U1918 (.A1(W624), .A2(W924), .ZN(W1918));
	INVX1 U1923 (.I(O173), .ZN(W1923));
	NANDX1 U1927 (.A1(W747), .A2(I1341), .ZN(W1927));
	NOR2X1 U1928 (.A1(I4493), .A2(W1168), .ZN(O3));
	NOR2X1 U1930 (.A1(W575), .A2(W888), .ZN(W1930));
	NANDX1 U1931 (.A1(I3388), .A2(W1289), .ZN(W1931));
	INVX1 U1932 (.I(W991), .ZN(W1932));
	NOR2X1 U1934 (.A1(W1458), .A2(I2896), .ZN(W1934));
	NANDX1 U1936 (.A1(W676), .A2(W498), .ZN(O498));
	INVX1 U1939 (.I(W1610), .ZN(O436));
	NANDX1 U1942 (.A1(I2355), .A2(I4805), .ZN(W1942));
	INVX1 U1944 (.I(W604), .ZN(W1944));
	NOR2X1 U1946 (.A1(W1179), .A2(W1434), .ZN(W1946));
	NOR2X1 U1948 (.A1(W637), .A2(I3335), .ZN(W1948));
	NANDX1 U1951 (.A1(I2566), .A2(I244), .ZN(W1951));
	INVX1 U1955 (.I(W1489), .ZN(O450));
	NANDX1 U1956 (.A1(W1799), .A2(I3532), .ZN(W1956));
	INVX1 U1959 (.I(W1185), .ZN(W1959));
	INVX1 U1960 (.I(W1655), .ZN(W1960));
	NOR2X1 U1961 (.A1(I2421), .A2(I3095), .ZN(W1961));
	NANDX1 U1963 (.A1(I903), .A2(W619), .ZN(W1963));
	NANDX1 U1966 (.A1(W1374), .A2(W45), .ZN(W1966));
	NOR2X1 U1970 (.A1(W664), .A2(I926), .ZN(W1970));
	NOR2X1 U1976 (.A1(W1679), .A2(W1470), .ZN(W1976));
	NOR2X1 U1980 (.A1(I4166), .A2(I1983), .ZN(W1980));
	NOR2X1 U1981 (.A1(I4885), .A2(W1801), .ZN(W1981));
	INVX1 U1982 (.I(I396), .ZN(W1982));
	NANDX1 U1991 (.A1(W987), .A2(I1130), .ZN(O43));
	NOR2X1 U1998 (.A1(W1981), .A2(I2060), .ZN(W1998));
	INVX1 U2005 (.I(W8), .ZN(W2005));
	INVX1 U2007 (.I(I2630), .ZN(W2007));
	NOR2X1 U2010 (.A1(I3352), .A2(I1558), .ZN(W2010));
	INVX1 U2012 (.I(W1604), .ZN(W2012));
	INVX1 U2013 (.I(I1287), .ZN(O239));
	NANDX1 U2018 (.A1(W409), .A2(I1287), .ZN(W2018));
	NANDX1 U2019 (.A1(I3787), .A2(W1680), .ZN(W2019));
	NOR2X1 U2031 (.A1(I4570), .A2(I594), .ZN(W2031));
	NANDX1 U2035 (.A1(O165), .A2(W85), .ZN(W2035));
	INVX1 U2040 (.I(I1943), .ZN(W2040));
	NANDX1 U2041 (.A1(I111), .A2(W626), .ZN(O469));
	INVX1 U2045 (.I(W108), .ZN(W2045));
	NOR2X1 U2047 (.A1(I3351), .A2(I2653), .ZN(W2047));
	NANDX1 U2048 (.A1(W1242), .A2(I2134), .ZN(W2048));
	NANDX1 U2050 (.A1(W1345), .A2(I2346), .ZN(W2050));
	INVX1 U2053 (.I(I4297), .ZN(W2053));
	NANDX1 U2057 (.A1(I1297), .A2(W1284), .ZN(W2057));
	NOR2X1 U2061 (.A1(I1528), .A2(I4584), .ZN(W2061));
	NANDX1 U2066 (.A1(W22), .A2(W1942), .ZN(W2066));
	NOR2X1 U2069 (.A1(W1661), .A2(I1506), .ZN(O314));
	NANDX1 U2070 (.A1(W838), .A2(W1069), .ZN(W2070));
	NOR2X1 U2072 (.A1(I2859), .A2(I1341), .ZN(W2072));
	NANDX1 U2080 (.A1(I4600), .A2(W150), .ZN(W2080));
	NOR2X1 U2082 (.A1(I4227), .A2(I434), .ZN(O380));
	NANDX1 U2083 (.A1(W800), .A2(I1565), .ZN(W2083));
	INVX1 U2085 (.I(W854), .ZN(W2085));
	NANDX1 U2087 (.A1(W1490), .A2(I541), .ZN(W2087));
	NANDX1 U2088 (.A1(W639), .A2(I2972), .ZN(O306));
	NANDX1 U2093 (.A1(W1357), .A2(I960), .ZN(W2093));
	INVX1 U2099 (.I(W1719), .ZN(W2099));
	NOR2X1 U2101 (.A1(I2644), .A2(W864), .ZN(W2101));
	NANDX1 U2103 (.A1(I2976), .A2(W1593), .ZN(W2103));
	NANDX1 U2115 (.A1(I1578), .A2(W1301), .ZN(W2115));
	NANDX1 U2121 (.A1(W1158), .A2(W952), .ZN(W2121));
	NOR2X1 U2127 (.A1(W896), .A2(I2645), .ZN(O257));
	NOR2X1 U2131 (.A1(W515), .A2(I2474), .ZN(W2131));
	NOR2X1 U2136 (.A1(W625), .A2(W1430), .ZN(W2136));
	NOR2X1 U2138 (.A1(I2842), .A2(W297), .ZN(W2138));
	NANDX1 U2141 (.A1(I480), .A2(I4042), .ZN(O93));
	NOR2X1 U2142 (.A1(I4327), .A2(W697), .ZN(W2142));
	NANDX1 U2144 (.A1(I3672), .A2(I3915), .ZN(W2144));
	NANDX1 U2146 (.A1(I4910), .A2(I2338), .ZN(W2146));
	NOR2X1 U2147 (.A1(W1574), .A2(W1037), .ZN(W2147));
	INVX1 U2151 (.I(W1091), .ZN(W2151));
	NANDX1 U2154 (.A1(I58), .A2(W458), .ZN(W2154));
	NANDX1 U2160 (.A1(W1420), .A2(W74), .ZN(O42));
	NANDX1 U2169 (.A1(W1744), .A2(I605), .ZN(W2169));
	NANDX1 U2171 (.A1(O314), .A2(I1894), .ZN(W2171));
	INVX1 U2178 (.I(I4466), .ZN(W2178));
	NANDX1 U2183 (.A1(W1028), .A2(I579), .ZN(W2183));
	NANDX1 U2184 (.A1(W1273), .A2(I1373), .ZN(W2184));
	NANDX1 U2188 (.A1(I3114), .A2(W556), .ZN(W2188));
	NANDX1 U2189 (.A1(W1066), .A2(W1721), .ZN(W2189));
	NOR2X1 U2194 (.A1(I4020), .A2(W2007), .ZN(W2194));
	NANDX1 U2196 (.A1(W196), .A2(I4063), .ZN(W2196));
	NANDX1 U2203 (.A1(W649), .A2(O420), .ZN(W2203));
	NOR2X1 U2206 (.A1(W728), .A2(I1535), .ZN(O29));
	NANDX1 U2208 (.A1(I3883), .A2(I2438), .ZN(W2208));
	NOR2X1 U2212 (.A1(W249), .A2(W2188), .ZN(W2212));
	INVX1 U2216 (.I(I3847), .ZN(W2216));
	NOR2X1 U2223 (.A1(W0), .A2(W541), .ZN(W2223));
	NANDX1 U2225 (.A1(I3623), .A2(W1272), .ZN(W2225));
	NANDX1 U2230 (.A1(I2704), .A2(W1462), .ZN(W2230));
	INVX1 U2235 (.I(W2083), .ZN(W2235));
	INVX1 U2237 (.I(W2212), .ZN(W2237));
	INVX1 U2239 (.I(I1535), .ZN(W2239));
	INVX1 U2247 (.I(O283), .ZN(W2247));
	NOR2X1 U2254 (.A1(I2929), .A2(I3816), .ZN(W2254));
	NANDX1 U2255 (.A1(O482), .A2(W426), .ZN(O76));
	NANDX1 U2259 (.A1(W593), .A2(W1040), .ZN(W2259));
	INVX1 U2262 (.I(I1890), .ZN(O358));
	NANDX1 U2264 (.A1(W1895), .A2(W649), .ZN(W2264));
	NOR2X1 U2266 (.A1(W826), .A2(I545), .ZN(W2266));
	NOR2X1 U2267 (.A1(W1890), .A2(W2005), .ZN(W2267));
	NOR2X1 U2277 (.A1(W2099), .A2(I4215), .ZN(W2277));
	NOR2X1 U2278 (.A1(W1242), .A2(I940), .ZN(W2278));
	NANDX1 U2281 (.A1(I2278), .A2(W157), .ZN(O55));
	NANDX1 U2282 (.A1(I929), .A2(W1373), .ZN(W2282));
	NOR2X1 U2283 (.A1(I3936), .A2(W2178), .ZN(W2283));
	NOR2X1 U2290 (.A1(I615), .A2(W600), .ZN(O456));
	NANDX1 U2293 (.A1(I4307), .A2(I3268), .ZN(W2293));
	NOR2X1 U2294 (.A1(I3448), .A2(W2277), .ZN(W2294));
	INVX1 U2296 (.I(I4603), .ZN(W2296));
	INVX1 U2297 (.I(W1747), .ZN(W2297));
	NANDX1 U2298 (.A1(I440), .A2(I114), .ZN(W2298));
	INVX1 U2302 (.I(W1736), .ZN(W2302));
	NANDX1 U2311 (.A1(I4328), .A2(I643), .ZN(O123));
	INVX1 U2313 (.I(I1724), .ZN(W2313));
	NOR2X1 U2316 (.A1(W1225), .A2(I675), .ZN(W2316));
	NOR2X1 U2320 (.A1(W1237), .A2(W18), .ZN(W2320));
	INVX1 U2321 (.I(W2053), .ZN(W2321));
	INVX1 U2327 (.I(W2066), .ZN(W2327));
	INVX1 U2329 (.I(W1813), .ZN(W2329));
	NANDX1 U2331 (.A1(I3816), .A2(W1275), .ZN(W2331));
	NOR2X1 U2333 (.A1(I1132), .A2(W1405), .ZN(O67));
	INVX1 U2335 (.I(W617), .ZN(W2335));
	NANDX1 U2339 (.A1(I4061), .A2(W869), .ZN(W2339));
	NOR2X1 U2340 (.A1(W1797), .A2(W1690), .ZN(W2340));
	NOR2X1 U2341 (.A1(I40), .A2(I3444), .ZN(W2341));
	NANDX1 U2343 (.A1(I4658), .A2(W1382), .ZN(W2343));
	INVX1 U2346 (.I(W2343), .ZN(W2346));
	INVX1 U2349 (.I(W428), .ZN(W2349));
	INVX1 U2354 (.I(W1527), .ZN(W2354));
	NANDX1 U2362 (.A1(W1120), .A2(W220), .ZN(W2362));
	NANDX1 U2375 (.A1(I4719), .A2(W1372), .ZN(W2375));
	NANDX1 U2382 (.A1(W2169), .A2(I4462), .ZN(W2382));
	INVX1 U2386 (.I(W1960), .ZN(W2386));
	INVX1 U2387 (.I(I937), .ZN(W2387));
	NANDX1 U2388 (.A1(W1585), .A2(I963), .ZN(O117));
	NOR2X1 U2389 (.A1(I1291), .A2(I4753), .ZN(W2389));
	NANDX1 U2392 (.A1(I3408), .A2(I1314), .ZN(W2392));
	NOR2X1 U2394 (.A1(O408), .A2(I2254), .ZN(W2394));
	NANDX1 U2398 (.A1(I380), .A2(I2882), .ZN(W2398));
	NOR2X1 U2400 (.A1(W10), .A2(W788), .ZN(W2400));
	NANDX1 U2403 (.A1(W2239), .A2(W157), .ZN(W2403));
	INVX1 U2408 (.I(W2099), .ZN(W2408));
	INVX1 U2410 (.I(I1314), .ZN(W2410));
	NOR2X1 U2411 (.A1(I347), .A2(I3018), .ZN(W2411));
	NANDX1 U2413 (.A1(O42), .A2(I3999), .ZN(W2413));
	INVX1 U2416 (.I(W2392), .ZN(W2416));
	NOR2X1 U2418 (.A1(I2657), .A2(I974), .ZN(W2418));
	INVX1 U2422 (.I(W909), .ZN(W2422));
	NANDX1 U2427 (.A1(I4611), .A2(W646), .ZN(W2427));
	INVX1 U2433 (.I(I2491), .ZN(O292));
	INVX1 U2434 (.I(W992), .ZN(O352));
	INVX1 U2436 (.I(O459), .ZN(W2436));
	NANDX1 U2438 (.A1(W122), .A2(I2062), .ZN(W2438));
	INVX1 U2439 (.I(I538), .ZN(W2439));
	INVX1 U2441 (.I(I1287), .ZN(W2441));
	NOR2X1 U2453 (.A1(W1558), .A2(W983), .ZN(W2453));
	NOR2X1 U2455 (.A1(I3219), .A2(I459), .ZN(W2455));
	NOR2X1 U2456 (.A1(W2035), .A2(I1498), .ZN(W2456));
	INVX1 U2465 (.I(I4257), .ZN(W2465));
	NANDX1 U2468 (.A1(W873), .A2(W1966), .ZN(W2468));
	NOR2X1 U2472 (.A1(W424), .A2(I4234), .ZN(W2472));
	NOR2X1 U2475 (.A1(W2189), .A2(I1615), .ZN(O148));
	NOR2X1 U2476 (.A1(W2394), .A2(W1345), .ZN(W2476));
	NANDX1 U2480 (.A1(I3381), .A2(W1509), .ZN(W2480));
	INVX1 U2483 (.I(W1725), .ZN(W2483));
	NANDX1 U2487 (.A1(I2974), .A2(W2320), .ZN(W2487));
	NANDX1 U2488 (.A1(W451), .A2(I4259), .ZN(W2488));
	NANDX1 U2489 (.A1(W1834), .A2(I2854), .ZN(W2489));
	NOR2X1 U2493 (.A1(I2731), .A2(I447), .ZN(W2493));
	INVX1 U2497 (.I(W2278), .ZN(W2497));
	NOR2X1 U2498 (.A1(W1503), .A2(I4293), .ZN(W2498));
	NOR2X1 U2507 (.A1(I2797), .A2(I2605), .ZN(W2507));
	NOR2X1 U2513 (.A1(W1868), .A2(W345), .ZN(W2513));
	NANDX1 U2514 (.A1(I4276), .A2(I1647), .ZN(W2514));
	NANDX1 U2524 (.A1(I1874), .A2(W205), .ZN(O189));
	NOR2X1 U2525 (.A1(O267), .A2(I748), .ZN(W2525));
	NOR2X1 U2528 (.A1(O192), .A2(W1732), .ZN(W2528));
	NOR2X1 U2547 (.A1(I3611), .A2(W2441), .ZN(W2547));
	NANDX1 U2549 (.A1(W2297), .A2(W2259), .ZN(O194));
	NOR2X1 U2552 (.A1(W1275), .A2(W783), .ZN(W2552));
	NANDX1 U2555 (.A1(I2046), .A2(W1930), .ZN(W2555));
	NOR2X1 U2561 (.A1(W1285), .A2(W2057), .ZN(W2561));
	INVX1 U2564 (.I(W1158), .ZN(O34));
	NANDX1 U2573 (.A1(I1179), .A2(W2410), .ZN(W2573));
	NANDX1 U2577 (.A1(W459), .A2(W1158), .ZN(W2577));
	NOR2X1 U2579 (.A1(W497), .A2(W959), .ZN(W2579));
	NOR2X1 U2584 (.A1(O42), .A2(O194), .ZN(W2584));
	NANDX1 U2587 (.A1(I3965), .A2(I2868), .ZN(W2587));
	NANDX1 U2589 (.A1(I630), .A2(I2962), .ZN(W2589));
	INVX1 U2598 (.I(I1391), .ZN(W2598));
	INVX1 U2604 (.I(I570), .ZN(W2604));
	INVX1 U2608 (.I(W1558), .ZN(O159));
	INVX1 U2613 (.I(W1693), .ZN(O238));
	NOR2X1 U2615 (.A1(I3928), .A2(I392), .ZN(O177));
	NANDX1 U2620 (.A1(I4135), .A2(W1341), .ZN(W2620));
	NOR2X1 U2622 (.A1(W1770), .A2(W630), .ZN(W2622));
	NOR2X1 U2626 (.A1(I3176), .A2(I2334), .ZN(O94));
	NANDX1 U2627 (.A1(W519), .A2(W1998), .ZN(W2627));
	INVX1 U2628 (.I(I3421), .ZN(W2628));
	NOR2X1 U2630 (.A1(W1044), .A2(I542), .ZN(W2630));
	INVX1 U2634 (.I(I4384), .ZN(W2634));
	NOR2X1 U2637 (.A1(I4160), .A2(I2434), .ZN(W2637));
	NOR2X1 U2648 (.A1(W2254), .A2(I3436), .ZN(W2648));
	NOR2X1 U2650 (.A1(I3984), .A2(W1430), .ZN(W2650));
	NOR2X1 U2653 (.A1(W35), .A2(W2403), .ZN(W2653));
	INVX1 U2663 (.I(W1568), .ZN(O155));
	NOR2X1 U2668 (.A1(I3930), .A2(W2099), .ZN(W2668));
	NOR2X1 U2670 (.A1(W771), .A2(I4703), .ZN(W2670));
	NANDX1 U2671 (.A1(W1188), .A2(I3543), .ZN(W2671));
	INVX1 U2676 (.I(W336), .ZN(W2676));
	NOR2X1 U2677 (.A1(W1096), .A2(W1795), .ZN(O339));
	INVX1 U2678 (.I(I4949), .ZN(O99));
	NOR2X1 U2682 (.A1(I4686), .A2(W1113), .ZN(W2682));
	NANDX1 U2683 (.A1(I14), .A2(I3394), .ZN(W2683));
	NANDX1 U2689 (.A1(W1624), .A2(I5), .ZN(W2689));
	NOR2X1 U2690 (.A1(I4831), .A2(I1913), .ZN(W2690));
	NANDX1 U2691 (.A1(I2238), .A2(W2398), .ZN(W2691));
	INVX1 U2692 (.I(I1292), .ZN(W2692));
	NOR2X1 U2696 (.A1(I2889), .A2(W2339), .ZN(W2696));
	INVX1 U2697 (.I(I4388), .ZN(W2697));
	NANDX1 U2699 (.A1(O21), .A2(W1874), .ZN(O153));
	NOR2X1 U2707 (.A1(I1541), .A2(I2408), .ZN(O434));
	INVX1 U2713 (.I(W471), .ZN(W2713));
	NANDX1 U2718 (.A1(W1319), .A2(W1850), .ZN(W2718));
	NANDX1 U2723 (.A1(I672), .A2(I1583), .ZN(W2723));
	NANDX1 U2725 (.A1(I1838), .A2(W2136), .ZN(W2725));
	INVX1 U2727 (.I(W1802), .ZN(W2727));
	NOR2X1 U2745 (.A1(I2880), .A2(W432), .ZN(W2745));
	INVX1 U2748 (.I(I1403), .ZN(O365));
	INVX1 U2753 (.I(W357), .ZN(W2753));
	INVX1 U2754 (.I(I4983), .ZN(W2754));
	NOR2X1 U2757 (.A1(W223), .A2(O267), .ZN(W2757));
	INVX1 U2758 (.I(W1910), .ZN(W2758));
	NOR2X1 U2764 (.A1(W1410), .A2(I3322), .ZN(W2764));
	NANDX1 U2771 (.A1(I3257), .A2(W458), .ZN(W2771));
	NOR2X1 U2772 (.A1(W119), .A2(W2223), .ZN(O134));
	NOR2X1 U2773 (.A1(W811), .A2(I4247), .ZN(O291));
	NOR2X1 U2775 (.A1(W224), .A2(I4597), .ZN(W2775));
	NANDX1 U2776 (.A1(W481), .A2(W2320), .ZN(O293));
	INVX1 U2783 (.I(I1274), .ZN(W2783));
	NOR2X1 U2786 (.A1(W1517), .A2(W788), .ZN(W2786));
	NOR2X1 U2789 (.A1(I4254), .A2(I4489), .ZN(W2789));
	INVX1 U2792 (.I(W1604), .ZN(W2792));
	NOR2X1 U2798 (.A1(I1535), .A2(W1815), .ZN(W2798));
	INVX1 U2803 (.I(W57), .ZN(W2803));
	NANDX1 U2806 (.A1(I863), .A2(I2094), .ZN(W2806));
	NOR2X1 U2812 (.A1(W2048), .A2(W988), .ZN(O312));
	NANDX1 U2818 (.A1(W2682), .A2(I919), .ZN(W2818));
	NANDX1 U2819 (.A1(I1608), .A2(I3688), .ZN(O454));
	NOR2X1 U2820 (.A1(W450), .A2(W1389), .ZN(O116));
	NANDX1 U2828 (.A1(W1357), .A2(I2859), .ZN(W2828));
	NANDX1 U2831 (.A1(I571), .A2(W125), .ZN(W2831));
	INVX1 U2835 (.I(W2313), .ZN(W2835));
	NOR2X1 U2837 (.A1(W2528), .A2(W2154), .ZN(W2837));
	NANDX1 U2842 (.A1(I2271), .A2(W2483), .ZN(W2842));
	NOR2X1 U2850 (.A1(W2453), .A2(W2386), .ZN(O415));
	NANDX1 U2852 (.A1(W1656), .A2(I59), .ZN(O274));
	NOR2X1 U2860 (.A1(W1915), .A2(W691), .ZN(O355));
	NOR2X1 U2864 (.A1(W229), .A2(W499), .ZN(W2864));
	NANDX1 U2872 (.A1(W1976), .A2(W2514), .ZN(O130));
	NOR2X1 U2880 (.A1(W1698), .A2(W2628), .ZN(O483));
	NOR2X1 U2881 (.A1(W419), .A2(I2588), .ZN(W2881));
	INVX1 U2889 (.I(O79), .ZN(W2889));
	NOR2X1 U2893 (.A1(W1247), .A2(W1400), .ZN(O199));
	NANDX1 U2894 (.A1(I1684), .A2(W487), .ZN(O139));
	INVX1 U2903 (.I(I2815), .ZN(W2903));
	NANDX1 U2910 (.A1(W1274), .A2(I4385), .ZN(W2910));
	NANDX1 U2926 (.A1(I857), .A2(W370), .ZN(O7));
	NOR2X1 U2928 (.A1(W2196), .A2(W1886), .ZN(W2928));
	INVX1 U2933 (.I(W430), .ZN(W2933));
	NOR2X1 U2936 (.A1(W1218), .A2(I2762), .ZN(O154));
	INVX1 U2937 (.I(W1363), .ZN(W2937));
	NANDX1 U2940 (.A1(W2622), .A2(I863), .ZN(O279));
	INVX1 U2949 (.I(W2648), .ZN(O263));
	NOR2X1 U2955 (.A1(I1185), .A2(W1742), .ZN(W2955));
	NANDX1 U2957 (.A1(W2389), .A2(I2926), .ZN(W2957));
	INVX1 U2958 (.I(W2346), .ZN(W2958));
	NANDX1 U2964 (.A1(W1948), .A2(W137), .ZN(W2964));
	NOR2X1 U2973 (.A1(I516), .A2(W1495), .ZN(W2973));
	NANDX1 U2974 (.A1(W195), .A2(W33), .ZN(W2974));
	NANDX1 U2979 (.A1(W2696), .A2(O99), .ZN(W2979));
	INVX1 U2984 (.I(W2282), .ZN(W2984));
	NOR2X1 U2987 (.A1(W1956), .A2(W1069), .ZN(W2987));
	NANDX1 U3002 (.A1(W2676), .A2(I107), .ZN(W3002));
	NANDX1 U3005 (.A1(I2037), .A2(W273), .ZN(W3005));
	NANDX1 U3013 (.A1(W807), .A2(W1216), .ZN(W3013));
	INVX1 U3014 (.I(W1931), .ZN(W3014));
	NOR2X1 U3021 (.A1(W2203), .A2(W1932), .ZN(W3021));
	INVX1 U3023 (.I(W92), .ZN(W3023));
	NOR2X1 U3032 (.A1(I2247), .A2(W2294), .ZN(W3032));
	NANDX1 U3035 (.A1(W3013), .A2(I1607), .ZN(O479));
	NOR2X1 U3036 (.A1(W2468), .A2(I1729), .ZN(W3036));
	NOR2X1 U3037 (.A1(W1185), .A2(W2555), .ZN(W3037));
	INVX1 U3052 (.I(I2365), .ZN(W3052));
	INVX1 U3053 (.I(I4405), .ZN(W3053));
	NOR2X1 U3054 (.A1(W2144), .A2(I4636), .ZN(O419));
	INVX1 U3066 (.I(W2061), .ZN(W3066));
	NOR2X1 U3071 (.A1(I601), .A2(I393), .ZN(O62));
	NANDX1 U3072 (.A1(W1946), .A2(I4771), .ZN(W3072));
	NOR2X1 U3075 (.A1(I2989), .A2(W899), .ZN(W3075));
	INVX1 U3082 (.I(I3582), .ZN(O19));
	NOR2X1 U3083 (.A1(I1478), .A2(W2493), .ZN(W3083));
	NANDX1 U3084 (.A1(W1329), .A2(I2445), .ZN(W3084));
	INVX1 U3089 (.I(W1537), .ZN(W3089));
	NANDX1 U3090 (.A1(W2230), .A2(I158), .ZN(W3090));
	INVX1 U3098 (.I(W1592), .ZN(O407));
	NOR2X1 U3099 (.A1(W775), .A2(W1747), .ZN(W3099));
	NOR2X1 U3102 (.A1(I1797), .A2(W1037), .ZN(O286));
	NOR2X1 U3104 (.A1(I2196), .A2(W904), .ZN(W3104));
	INVX1 U3105 (.I(W2955), .ZN(W3105));
	NANDX1 U3110 (.A1(I4102), .A2(O460), .ZN(W3110));
	INVX1 U3126 (.I(I566), .ZN(W3126));
	NOR2X1 U3127 (.A1(I4534), .A2(W2973), .ZN(W3127));
	NANDX1 U3132 (.A1(W2828), .A2(I99), .ZN(W3132));
	NANDX1 U3137 (.A1(I4361), .A2(W1960), .ZN(W3137));
	INVX1 U3138 (.I(W2386), .ZN(W3138));
	NOR2X1 U3139 (.A1(I1919), .A2(W1189), .ZN(O303));
	INVX1 U3141 (.I(W408), .ZN(W3141));
	NANDX1 U3144 (.A1(W784), .A2(W848), .ZN(W3144));
	NANDX1 U3156 (.A1(W189), .A2(W1214), .ZN(O401));
	NOR2X1 U3159 (.A1(W2979), .A2(I1767), .ZN(W3159));
	NOR2X1 U3164 (.A1(I2710), .A2(W1064), .ZN(W3164));
	NANDX1 U3176 (.A1(I4772), .A2(W2653), .ZN(W3176));
	NOR2X1 U3185 (.A1(W1927), .A2(W1961), .ZN(W3185));
	INVX1 U3191 (.I(W418), .ZN(O10));
	NOR2X1 U3192 (.A1(I4104), .A2(I1536), .ZN(W3192));
	NANDX1 U3198 (.A1(W161), .A2(W1477), .ZN(O384));
	NOR2X1 U3200 (.A1(I3769), .A2(W837), .ZN(O453));
	NOR2X1 U3203 (.A1(W856), .A2(I485), .ZN(W3203));
	NANDX1 U3205 (.A1(W1688), .A2(W88), .ZN(W3205));
	NANDX1 U3215 (.A1(W1736), .A2(W2670), .ZN(W3215));
	NANDX1 U3216 (.A1(W2422), .A2(I3747), .ZN(W3216));
	INVX1 U3221 (.I(I3971), .ZN(O373));
	INVX1 U3226 (.I(W2668), .ZN(W3226));
	INVX1 U3227 (.I(W1761), .ZN(W3227));
	NANDX1 U3228 (.A1(O293), .A2(I2653), .ZN(O13));
	NOR2X1 U3229 (.A1(W2783), .A2(I4185), .ZN(W3229));
	INVX1 U3237 (.I(I3193), .ZN(W3237));
	INVX1 U3246 (.I(W25), .ZN(W3246));
	NANDX1 U3247 (.A1(W3176), .A2(W405), .ZN(W3247));
	NANDX1 U3250 (.A1(W1982), .A2(O333), .ZN(W3250));
	INVX1 U3255 (.I(W2410), .ZN(O202));
	NANDX1 U3261 (.A1(I4033), .A2(I619), .ZN(W3261));
	INVX1 U3262 (.I(I2610), .ZN(O497));
	NOR2X1 U3265 (.A1(I1872), .A2(W2723), .ZN(W3265));
	NANDX1 U3269 (.A1(W3005), .A2(W3141), .ZN(O171));
	NOR2X1 U3271 (.A1(W878), .A2(W2507), .ZN(W3271));
	NOR2X1 U3278 (.A1(I701), .A2(W2050), .ZN(W3278));
	INVX1 U3279 (.I(W1474), .ZN(O426));
	NOR2X1 U3282 (.A1(W2598), .A2(I546), .ZN(W3282));
	NANDX1 U3288 (.A1(W2142), .A2(W693), .ZN(W3288));
	NANDX1 U3289 (.A1(I594), .A2(I1795), .ZN(W3289));
	NOR2X1 U3298 (.A1(I4141), .A2(I3333), .ZN(W3298));
	NOR2X1 U3301 (.A1(I3887), .A2(I3965), .ZN(W3301));
	NOR2X1 U3302 (.A1(I4337), .A2(I1880), .ZN(W3302));
	INVX1 U3304 (.I(W528), .ZN(O32));
	INVX1 U3307 (.I(W463), .ZN(O325));
	NOR2X1 U3314 (.A1(O456), .A2(O114), .ZN(O206));
	NANDX1 U3317 (.A1(W2354), .A2(W1370), .ZN(W3317));
	NOR2X1 U3318 (.A1(W1737), .A2(I1012), .ZN(W3318));
	INVX1 U3333 (.I(W1473), .ZN(W3333));
	NOR2X1 U3344 (.A1(I3028), .A2(I4082), .ZN(W3344));
	NOR2X1 U3352 (.A1(W1233), .A2(I1863), .ZN(W3352));
	NOR2X1 U3363 (.A1(W534), .A2(W2436), .ZN(W3363));
	NANDX1 U3368 (.A1(W2266), .A2(I3367), .ZN(W3368));
	NANDX1 U3376 (.A1(W12), .A2(W2283), .ZN(W3376));
	NANDX1 U3380 (.A1(I3750), .A2(W2340), .ZN(W3380));
	NOR2X1 U3381 (.A1(W21), .A2(W1415), .ZN(W3381));
	NOR2X1 U3394 (.A1(W787), .A2(W1344), .ZN(O127));
	INVX1 U3396 (.I(I1914), .ZN(O108));
	NANDX1 U3400 (.A1(W3261), .A2(W568), .ZN(W3400));
	INVX1 U3401 (.I(I4216), .ZN(O271));
	INVX1 U3403 (.I(I1142), .ZN(O226));
	INVX1 U3405 (.I(W2488), .ZN(W3405));
	NOR2X1 U3430 (.A1(I4118), .A2(O13), .ZN(W3430));
	INVX1 U3435 (.I(W640), .ZN(W3435));
	INVX1 U3437 (.I(W1469), .ZN(O376));
	NOR2X1 U3441 (.A1(W3075), .A2(W3014), .ZN(W3441));
	NANDX1 U3443 (.A1(W2831), .A2(W2650), .ZN(O477));
	INVX1 U3445 (.I(W2045), .ZN(W3445));
	INVX1 U3448 (.I(I3957), .ZN(W3448));
	NOR2X1 U3449 (.A1(I3330), .A2(W1948), .ZN(W3449));
	NANDX1 U3450 (.A1(W117), .A2(W2713), .ZN(W3450));
	NOR2X1 U3452 (.A1(W2403), .A2(I2201), .ZN(W3452));
	NOR2X1 U3453 (.A1(O189), .A2(W3449), .ZN(W3453));
	INVX1 U3455 (.I(W176), .ZN(O243));
	INVX1 U3457 (.I(W564), .ZN(W3457));
	INVX1 U3464 (.I(W914), .ZN(W3464));
	NANDX1 U3478 (.A1(I3610), .A2(W3452), .ZN(O351));
	INVX1 U3481 (.I(W1863), .ZN(W3481));
	INVX1 U3495 (.I(O293), .ZN(W3495));
	NOR2X1 U3497 (.A1(W1944), .A2(I3744), .ZN(W3497));
	NOR2X1 U3502 (.A1(I1404), .A2(I4169), .ZN(W3502));
	INVX1 U3506 (.I(I2025), .ZN(O133));
	NOR2X1 U3508 (.A1(I3408), .A2(W466), .ZN(O463));
	NOR2X1 U3510 (.A1(I1121), .A2(W1392), .ZN(O457));
	NOR2X1 U3520 (.A1(W2480), .A2(W548), .ZN(W3520));
	NOR2X1 U3528 (.A1(W1145), .A2(W766), .ZN(O362));
	NOR2X1 U3535 (.A1(I4991), .A2(O159), .ZN(W3535));
	NOR2X1 U3557 (.A1(I2809), .A2(W156), .ZN(O427));
	NOR2X1 U3560 (.A1(I1943), .A2(W1970), .ZN(W3560));
	NANDX1 U3562 (.A1(W2889), .A2(W2375), .ZN(W3562));
	NANDX1 U3565 (.A1(W1951), .A2(W3138), .ZN(W3565));
	NOR2X1 U3566 (.A1(W2881), .A2(W1823), .ZN(W3566));
	INVX1 U3572 (.I(I3652), .ZN(W3572));
	NANDX1 U3574 (.A1(I971), .A2(I4946), .ZN(O231));
	NOR2X1 U3584 (.A1(I3933), .A2(W625), .ZN(W3584));
	NOR2X1 U3591 (.A1(I1726), .A2(W1247), .ZN(W3591));
	NOR2X1 U3593 (.A1(I4185), .A2(I3279), .ZN(O216));
	INVX1 U3608 (.I(I220), .ZN(O418));
	INVX1 U3615 (.I(W1837), .ZN(O317));
	NANDX1 U3618 (.A1(W2465), .A2(W2552), .ZN(O371));
	NOR2X1 U3627 (.A1(I1364), .A2(W2472), .ZN(W3627));
	INVX1 U3629 (.I(W3090), .ZN(W3629));
	INVX1 U3632 (.I(W3089), .ZN(W3632));
	INVX1 U3633 (.I(W2264), .ZN(O449));
	NANDX1 U3636 (.A1(W1096), .A2(W2070), .ZN(W3636));
	NANDX1 U3637 (.A1(W1874), .A2(W2147), .ZN(W3637));
	INVX1 U3639 (.I(W991), .ZN(W3639));
	INVX1 U3645 (.I(I3276), .ZN(W3645));
	NANDX1 U3646 (.A1(W446), .A2(I3017), .ZN(W3646));
	NOR2X1 U3647 (.A1(W3144), .A2(I174), .ZN(W3647));
	NOR2X1 U3657 (.A1(W901), .A2(I3918), .ZN(W3657));
	INVX1 U3659 (.I(I3601), .ZN(W3659));
	NANDX1 U3660 (.A1(W1272), .A2(W3137), .ZN(O97));
	NOR2X1 U3663 (.A1(W2910), .A2(O4), .ZN(W3663));
	INVX1 U3664 (.I(W486), .ZN(W3664));
	NOR2X1 U3667 (.A1(I4211), .A2(I4212), .ZN(W3667));
	NANDX1 U3677 (.A1(O197), .A2(W1772), .ZN(W3677));
	INVX1 U3686 (.I(I4595), .ZN(W3686));
	INVX1 U3692 (.I(W1097), .ZN(O338));
	INVX1 U3698 (.I(W3636), .ZN(W3698));
	NANDX1 U3699 (.A1(W3298), .A2(W1502), .ZN(W3699));
	NANDX1 U3704 (.A1(W2798), .A2(I3658), .ZN(W3704));
	NANDX1 U3712 (.A1(W121), .A2(W3246), .ZN(W3712));
	NOR2X1 U3717 (.A1(W3481), .A2(O139), .ZN(W3717));
	NANDX1 U3718 (.A1(I3683), .A2(W3333), .ZN(W3718));
	INVX1 U3720 (.I(W2115), .ZN(O66));
	INVX1 U3723 (.I(I1480), .ZN(W3723));
	INVX1 U3734 (.I(I430), .ZN(W3734));
	NOR2X1 U3754 (.A1(W1718), .A2(I486), .ZN(O58));
	NOR2X1 U3762 (.A1(I701), .A2(I1767), .ZN(O285));
	INVX1 U3772 (.I(W3464), .ZN(O431));
	NANDX1 U3790 (.A1(W2296), .A2(W3445), .ZN(W3790));
	INVX1 U3799 (.I(W1476), .ZN(W3799));
	NOR2X1 U3809 (.A1(W260), .A2(I3093), .ZN(W3809));
	NOR2X1 U3810 (.A1(W1863), .A2(W1881), .ZN(W3810));
	NOR2X1 U3815 (.A1(W2031), .A2(W3072), .ZN(W3815));
	INVX1 U3816 (.I(W1944), .ZN(W3816));
	INVX1 U3826 (.I(W3717), .ZN(O25));
	NANDX1 U3827 (.A1(W3566), .A2(W3627), .ZN(W3827));
	NANDX1 U3829 (.A1(I2108), .A2(I4029), .ZN(O364));
	NOR2X1 U3833 (.A1(W1045), .A2(I4058), .ZN(W3833));
	INVX1 U3835 (.I(I3428), .ZN(O204));
	NANDX1 U3842 (.A1(W2764), .A2(W750), .ZN(W3842));
	NANDX1 U3843 (.A1(W2627), .A2(W2047), .ZN(W3843));
	NOR2X1 U3847 (.A1(W3445), .A2(W3497), .ZN(W3847));
	NANDX1 U3849 (.A1(W1408), .A2(W3560), .ZN(W3849));
	NANDX1 U3852 (.A1(I3485), .A2(I1140), .ZN(W3852));
	NOR2X1 U3859 (.A1(W3159), .A2(I4414), .ZN(W3859));
	NANDX1 U3860 (.A1(O231), .A2(W2335), .ZN(W3860));
	NANDX1 U3867 (.A1(I630), .A2(W2864), .ZN(W3867));
	NOR2X1 U3868 (.A1(I465), .A2(W2489), .ZN(W3868));
	NOR2X1 U3873 (.A1(W2727), .A2(O55), .ZN(W3873));
	INVX1 U3878 (.I(W2757), .ZN(W3878));
	NANDX1 U3893 (.A1(W1430), .A2(W1934), .ZN(O258));
	NANDX1 U3897 (.A1(W1770), .A2(O97), .ZN(W3897));
	INVX1 U3913 (.I(I4832), .ZN(W3913));
	INVX1 U3923 (.I(W3216), .ZN(W3923));
	NOR2X1 U3924 (.A1(W1351), .A2(W256), .ZN(W3924));
	NOR2X1 U3928 (.A1(I2456), .A2(W2584), .ZN(W3928));
	NOR2X1 U3937 (.A1(W1772), .A2(I4955), .ZN(W3937));
	INVX1 U3939 (.I(W652), .ZN(W3939));
	INVX1 U3942 (.I(W3572), .ZN(W3942));
	INVX1 U3949 (.I(W2745), .ZN(O256));
	NOR2X1 U3950 (.A1(W1469), .A2(O441), .ZN(W3950));
	INVX1 U3951 (.I(I3114), .ZN(O128));
	NOR2X1 U3953 (.A1(W1380), .A2(W1657), .ZN(W3953));
	NOR2X1 U3955 (.A1(W3686), .A2(W713), .ZN(W3955));
	NANDX1 U3958 (.A1(W3937), .A2(W414), .ZN(O255));
	NOR2X1 U3963 (.A1(W2468), .A2(I2575), .ZN(O368));
	NOR2X1 U3968 (.A1(W3368), .A2(W1178), .ZN(W3968));
	NANDX1 U3970 (.A1(W2093), .A2(W3924), .ZN(W3970));
	NANDX1 U3973 (.A1(W2121), .A2(I3986), .ZN(O318));
	NANDX1 U3974 (.A1(I1049), .A2(I1200), .ZN(W3974));
	INVX1 U3983 (.I(I2801), .ZN(W3983));
	INVX1 U3986 (.I(W3282), .ZN(W3986));
	NANDX1 U3991 (.A1(W3099), .A2(I3895), .ZN(W3991));
	NANDX1 U3993 (.A1(O449), .A2(W1874), .ZN(W3993));
	INVX1 U3994 (.I(W3698), .ZN(W3994));
	NANDX1 U3999 (.A1(W805), .A2(I4900), .ZN(W3999));
	NOR2X1 U4001 (.A1(W2138), .A2(W3192), .ZN(O200));
	INVX1 U4002 (.I(W3842), .ZN(O354));
	INVX1 U4004 (.I(I1550), .ZN(W4004));
	NOR2X1 U4017 (.A1(W908), .A2(W3712), .ZN(W4017));
	INVX1 U4033 (.I(W2171), .ZN(W4033));
	INVX1 U4035 (.I(W3535), .ZN(W4035));
	NOR2X1 U4063 (.A1(W2010), .A2(W2758), .ZN(W4063));
	NANDX1 U4065 (.A1(I1147), .A2(W2151), .ZN(W4065));
	INVX1 U4079 (.I(W3250), .ZN(W4079));
	INVX1 U4083 (.I(W2298), .ZN(W4083));
	INVX1 U4084 (.I(W2589), .ZN(W4084));
	NOR2X1 U4094 (.A1(I540), .A2(W3110), .ZN(O27));
	INVX1 U4097 (.I(W3913), .ZN(W4097));
	INVX1 U4112 (.I(I3127), .ZN(W4112));
	INVX1 U4113 (.I(W1293), .ZN(W4113));
	NANDX1 U4115 (.A1(W3226), .A2(W1998), .ZN(W4115));
	NANDX1 U4118 (.A1(W3860), .A2(W1697), .ZN(W4118));
	NANDX1 U4119 (.A1(I4026), .A2(I1179), .ZN(O212));
	NANDX1 U4121 (.A1(W8), .A2(W3363), .ZN(W4121));
	INVX1 U4123 (.I(W2321), .ZN(O35));
	NOR2X1 U4124 (.A1(W3704), .A2(I4669), .ZN(O104));
	INVX1 U4129 (.I(W276), .ZN(W4129));
	INVX1 U4131 (.I(I3401), .ZN(W4131));
	NOR2X1 U4135 (.A1(W2101), .A2(I2126), .ZN(O80));
	NOR2X1 U4138 (.A1(W3502), .A2(W1297), .ZN(W4138));
	NANDX1 U4139 (.A1(W3663), .A2(O74), .ZN(W4139));
	NANDX1 U4162 (.A1(I3441), .A2(I3991), .ZN(O356));
	INVX1 U4163 (.I(I4005), .ZN(W4163));
	NOR2X1 U4164 (.A1(I4850), .A2(W2455), .ZN(W4164));
	NANDX1 U4214 (.A1(I2344), .A2(I4118), .ZN(W4214));
	INVX1 U4229 (.I(I1518), .ZN(W4229));
	INVX1 U4237 (.I(W151), .ZN(O316));
	NOR2X1 U4259 (.A1(I2284), .A2(I1262), .ZN(W4259));
	NOR2X1 U4264 (.A1(I1300), .A2(W2671), .ZN(W4264));
	NOR2X1 U4267 (.A1(W1045), .A2(W884), .ZN(W4267));
	INVX1 U4271 (.I(W3809), .ZN(W4271));
	NANDX1 U4272 (.A1(I1256), .A2(I4106), .ZN(O277));
	NOR2X1 U4276 (.A1(W2235), .A2(W606), .ZN(O298));
	NANDX1 U4283 (.A1(W2933), .A2(W665), .ZN(W4283));
	INVX1 U4294 (.I(W426), .ZN(W4294));
	NOR2X1 U4296 (.A1(W3809), .A2(W1539), .ZN(W4296));
	INVX1 U4302 (.I(W2018), .ZN(W4302));
	NOR2X1 U4304 (.A1(I1654), .A2(W2690), .ZN(W4304));
	INVX1 U4305 (.I(W323), .ZN(W4305));
	INVX1 U4323 (.I(W2775), .ZN(W4323));
	NANDX1 U4325 (.A1(W686), .A2(W1433), .ZN(W4325));
	NANDX1 U4334 (.A1(W596), .A2(I3562), .ZN(W4334));
	NOR2X1 U4339 (.A1(W842), .A2(W2329), .ZN(O236));
	INVX1 U4347 (.I(W3448), .ZN(W4347));
	INVX1 U4357 (.I(I431), .ZN(W4357));
	NANDX1 U4367 (.A1(W964), .A2(W440), .ZN(W4367));
	NOR2X1 U4385 (.A1(W1320), .A2(I1690), .ZN(O402));
	INVX1 U4393 (.I(W4283), .ZN(O49));
	NANDX1 U4397 (.A1(W3464), .A2(W1154), .ZN(O143));
	INVX1 U4400 (.I(W3993), .ZN(O390));
	NANDX1 U4412 (.A1(O62), .A2(W3942), .ZN(W4412));
	NOR2X1 U4414 (.A1(W3053), .A2(I2319), .ZN(W4414));
	INVX1 U4421 (.I(W1779), .ZN(W4421));
	INVX1 U4423 (.I(W1396), .ZN(W4423));
	NANDX1 U4425 (.A1(W1769), .A2(W3827), .ZN(O115));
	NOR2X1 U4433 (.A1(W248), .A2(W4138), .ZN(W4433));
	INVX1 U4435 (.I(W4097), .ZN(W4435));
	NOR2X1 U4437 (.A1(W106), .A2(W2480), .ZN(O86));
	NOR2X1 U4438 (.A1(I3958), .A2(W2637), .ZN(W4438));
	NANDX1 U4440 (.A1(W4294), .A2(W2316), .ZN(W4440));
	NANDX1 U4441 (.A1(I1720), .A2(I758), .ZN(O39));
	INVX1 U4447 (.I(W3002), .ZN(O332));
	NOR2X1 U4449 (.A1(O394), .A2(W3066), .ZN(O217));
	NOR2X1 U4451 (.A1(I769), .A2(W1304), .ZN(W4451));
	INVX1 U4453 (.I(W196), .ZN(W4453));
	NANDX1 U4459 (.A1(I1154), .A2(I3801), .ZN(O471));
	NANDX1 U4466 (.A1(O463), .A2(W1633), .ZN(W4466));
	NANDX1 U4468 (.A1(O395), .A2(I2068), .ZN(W4468));
	NOR2X1 U4476 (.A1(W2266), .A2(W1140), .ZN(W4476));
	NANDX1 U4478 (.A1(W2087), .A2(W488), .ZN(W4478));
	NOR2X1 U4488 (.A1(I1932), .A2(W2842), .ZN(W4488));
	NANDX1 U4493 (.A1(I2970), .A2(W1589), .ZN(O51));
	NOR2X1 U4498 (.A1(W2903), .A2(W3632), .ZN(O46));
	NOR2X1 U4499 (.A1(W2382), .A2(I754), .ZN(W4499));
	NANDX1 U4505 (.A1(W1219), .A2(W3983), .ZN(O300));
	NOR2X1 U4508 (.A1(O183), .A2(W1401), .ZN(W4508));
	INVX1 U4511 (.I(I3351), .ZN(O272));
	NANDX1 U4516 (.A1(W1050), .A2(W4131), .ZN(W4516));
	INVX1 U4517 (.I(W4079), .ZN(W4517));
	INVX1 U4529 (.I(W980), .ZN(O210));
	NOR2X1 U4538 (.A1(W4302), .A2(W488), .ZN(O379));
	INVX1 U4552 (.I(W1328), .ZN(W4552));
	NANDX1 U4556 (.A1(W3986), .A2(W2438), .ZN(O363));
	NOR2X1 U4560 (.A1(W2771), .A2(W3271), .ZN(O472));
	NANDX1 U4572 (.A1(I4196), .A2(W3250), .ZN(W4572));
	NANDX1 U4573 (.A1(W1741), .A2(W4438), .ZN(W4573));
	INVX1 U4578 (.I(W112), .ZN(O391));
	NANDX1 U4597 (.A1(O115), .A2(W3203), .ZN(W4597));
	NANDX1 U4598 (.A1(W929), .A2(W2103), .ZN(W4598));
	NOR2X1 U4601 (.A1(W1540), .A2(W2835), .ZN(W4601));
	NANDX1 U4607 (.A1(W915), .A2(I3393), .ZN(W4607));
	INVX1 U4608 (.I(W2387), .ZN(W4608));
	NANDX1 U4619 (.A1(W1714), .A2(W2418), .ZN(W4619));
	NOR2X1 U4626 (.A1(W1571), .A2(W802), .ZN(W4626));
	INVX1 U4630 (.I(W577), .ZN(W4630));
	NANDX1 U4635 (.A1(W4451), .A2(W2573), .ZN(W4635));
	NOR2X1 U4638 (.A1(W4004), .A2(W4323), .ZN(W4638));
	INVX1 U4647 (.I(W3023), .ZN(O119));
	NOR2X1 U4651 (.A1(W1190), .A2(W120), .ZN(W4651));
	INVX1 U4654 (.I(I4112), .ZN(O220));
	NOR2X1 U4657 (.A1(I3241), .A2(W3847), .ZN(W4657));
	NANDX1 U4666 (.A1(W398), .A2(I894), .ZN(O430));
	NOR2X1 U4673 (.A1(W4635), .A2(W3734), .ZN(W4673));
	INVX1 U4688 (.I(O51), .ZN(W4688));
	NANDX1 U4697 (.A1(W3645), .A2(I561), .ZN(W4697));
	NANDX1 U4699 (.A1(W4516), .A2(W4433), .ZN(O280));
	INVX1 U4706 (.I(W729), .ZN(W4706));
	INVX1 U4721 (.I(O408), .ZN(O400));
	INVX1 U4726 (.I(I3653), .ZN(O490));
	NOR2X1 U4733 (.A1(I544), .A2(W4083), .ZN(O437));
	NANDX1 U4738 (.A1(W3302), .A2(W2964), .ZN(W4738));
	NOR2X1 U4754 (.A1(W960), .A2(I3222), .ZN(W4754));
	NOR2X1 U4794 (.A1(I562), .A2(W1386), .ZN(W4794));
	INVX1 U4799 (.I(W4115), .ZN(W4799));
	NOR2X1 U4812 (.A1(W3318), .A2(W3816), .ZN(O353));
	INVX1 U4818 (.I(W4347), .ZN(O476));
	NOR2X1 U4822 (.A1(W3718), .A2(I2812), .ZN(W4822));
	NOR2X1 U4824 (.A1(I3703), .A2(W3970), .ZN(W4824));
	NANDX1 U4825 (.A1(I2071), .A2(W4264), .ZN(O289));
	NOR2X1 U4828 (.A1(W3664), .A2(W2362), .ZN(W4828));
	NOR2X1 U4831 (.A1(W1019), .A2(I3388), .ZN(W4831));
	INVX1 U4859 (.I(W3205), .ZN(O221));
	NOR2X1 U4865 (.A1(W2525), .A2(O265), .ZN(W4865));
	NOR2X1 U4883 (.A1(W1470), .A2(W1048), .ZN(W4883));
	NANDX1 U4886 (.A1(W3520), .A2(W4259), .ZN(W4886));
	NANDX1 U4901 (.A1(W637), .A2(W159), .ZN(O248));
	NANDX1 U4909 (.A1(W2579), .A2(I3618), .ZN(W4909));
	NANDX1 U4911 (.A1(W1541), .A2(I3865), .ZN(O149));
	INVX1 U4919 (.I(W4084), .ZN(W4919));
	INVX1 U4920 (.I(W2341), .ZN(W4920));
	NOR2X1 U4923 (.A1(W2072), .A2(W1205), .ZN(O57));
	NANDX1 U4933 (.A1(O134), .A2(I4050), .ZN(O464));
	INVX1 U4938 (.I(O390), .ZN(W4938));
	NANDX1 U4947 (.A1(I1767), .A2(W3994), .ZN(W4947));
	NOR2X1 U4959 (.A1(O363), .A2(W1194), .ZN(W4959));
	NANDX1 U4962 (.A1(W764), .A2(W2634), .ZN(W4962));
	NOR2X1 U4965 (.A1(W1762), .A2(W3815), .ZN(W4965));
	NANDX1 U4966 (.A1(I1286), .A2(W731), .ZN(W4966));
	INVX1 U4974 (.I(W1234), .ZN(O488));
	INVX1 U4983 (.I(W4367), .ZN(O120));
	NANDX1 U4985 (.A1(I1482), .A2(I416), .ZN(W4985));
	INVX1 U4991 (.I(W284), .ZN(W4991));
	NANDX1 U4993 (.A1(O58), .A2(W3639), .ZN(W4993));
	NANDX1 U4994 (.A1(I54), .A2(W2184), .ZN(O84));
	INVX1 U5009 (.I(W1959), .ZN(W5009));
	NANDX1 U5013 (.A1(W2085), .A2(W1138), .ZN(W5013));
	NOR2X1 U5027 (.A1(W4630), .A2(I4860), .ZN(W5027));
	NANDX1 U5034 (.A1(W2561), .A2(W3849), .ZN(O275));
	NOR2X1 U5036 (.A1(W1718), .A2(I2595), .ZN(W5036));
	NANDX1 U5044 (.A1(I4325), .A2(W3867), .ZN(O466));
	NOR2X1 U5049 (.A1(W1536), .A2(O34), .ZN(W5049));
	NANDX1 U5054 (.A1(W1322), .A2(W3659), .ZN(W5054));
	NOR2X1 U5065 (.A1(W3974), .A2(W2577), .ZN(O309));
	INVX1 U5069 (.I(W1324), .ZN(W5069));
	INVX1 U5073 (.I(W4017), .ZN(W5073));
	INVX1 U5088 (.I(W4828), .ZN(W5088));
	NANDX1 U5099 (.A1(W36), .A2(O256), .ZN(W5099));
	NOR2X1 U5101 (.A1(W3132), .A2(I4292), .ZN(W5101));
	NANDX1 U5107 (.A1(W4962), .A2(I3783), .ZN(O480));
	NOR2X1 U5113 (.A1(W1405), .A2(W3450), .ZN(W5113));
	INVX1 U5116 (.I(W324), .ZN(O383));
	NANDX1 U5117 (.A1(W1439), .A2(W3999), .ZN(W5117));
	NANDX1 U5125 (.A1(W487), .A2(W607), .ZN(W5125));
	NOR2X1 U5146 (.A1(I2570), .A2(I2020), .ZN(O224));
	NANDX1 U5153 (.A1(I3344), .A2(W1192), .ZN(W5153));
	NANDX1 U5170 (.A1(I4180), .A2(W5049), .ZN(O105));
	NOR2X1 U5171 (.A1(W5027), .A2(W3381), .ZN(O52));
	INVX1 U5174 (.I(I332), .ZN(W5174));
	NANDX1 U5190 (.A1(W4113), .A2(W1372), .ZN(O294));
	INVX1 U5197 (.I(W3352), .ZN(W5197));
	INVX1 U5211 (.I(W3939), .ZN(W5211));
	NANDX1 U5218 (.A1(W2692), .A2(W3923), .ZN(O323));
	NOR2X1 U5229 (.A1(W2400), .A2(O130), .ZN(W5229));
	NANDX1 U5231 (.A1(W424), .A2(W476), .ZN(W5231));
	NANDX1 U5233 (.A1(W2803), .A2(I4627), .ZN(W5233));
	NOR2X1 U5235 (.A1(O161), .A2(I4363), .ZN(W5235));
	NANDX1 U5239 (.A1(I818), .A2(W1069), .ZN(O157));
	INVX1 U5241 (.I(I2219), .ZN(W5241));
	NOR2X1 U5251 (.A1(W5229), .A2(W2958), .ZN(O250));
	NOR2X1 U5276 (.A1(W4651), .A2(W2806), .ZN(W5276));
	NOR2X1 U5278 (.A1(W1039), .A2(W1304), .ZN(W5278));
	NANDX1 U5283 (.A1(W1301), .A2(I2072), .ZN(W5283));
	NOR2X1 U5284 (.A1(I3349), .A2(W1388), .ZN(O262));
	NOR2X1 U5302 (.A1(I3099), .A2(W4112), .ZN(O0));
	INVX1 U5306 (.I(W4626), .ZN(O372));
	NANDX1 U5324 (.A1(W882), .A2(W4688), .ZN(W5324));
	INVX1 U5327 (.I(W1387), .ZN(W5327));
	NANDX1 U5331 (.A1(W5069), .A2(W5278), .ZN(O168));
	NANDX1 U5332 (.A1(W3667), .A2(W3677), .ZN(O178));
	INVX1 U5333 (.I(W3647), .ZN(W5333));
	NOR2X1 U5334 (.A1(W445), .A2(W2439), .ZN(W5334));
	NANDX1 U5336 (.A1(W2691), .A2(W4638), .ZN(W5336));
	INVX1 U5338 (.I(W1561), .ZN(O121));
	NANDX1 U5347 (.A1(W4601), .A2(W5327), .ZN(O151));
	INVX1 U5356 (.I(I2561), .ZN(W5356));
	INVX1 U5360 (.I(I3236), .ZN(O14));
	NANDX1 U5363 (.A1(W3868), .A2(I1140), .ZN(W5363));
	NANDX1 U5372 (.A1(O176), .A2(W4478), .ZN(W5372));
	INVX1 U5373 (.I(I2694), .ZN(W5373));
	NANDX1 U5375 (.A1(W4697), .A2(O298), .ZN(W5375));
	INVX1 U5378 (.I(W265), .ZN(W5378));
	NOR2X1 U5382 (.A1(I579), .A2(W3441), .ZN(W5382));
	NANDX1 U5383 (.A1(W3790), .A2(I987), .ZN(O98));
	NANDX1 U5384 (.A1(W3584), .A2(W2587), .ZN(O92));
	INVX1 U5388 (.I(W3453), .ZN(W5388));
	INVX1 U5403 (.I(W1562), .ZN(W5403));
	NANDX1 U5404 (.A1(I777), .A2(W3572), .ZN(W5404));
	NOR2X1 U5405 (.A1(W4214), .A2(I4596), .ZN(W5405));
	NOR2X1 U5417 (.A1(W5276), .A2(W4453), .ZN(O190));
	NOR2X1 U5425 (.A1(W5231), .A2(W803), .ZN(O315));
	NOR2X1 U5426 (.A1(I2412), .A2(W1918), .ZN(W5426));
	NOR2X1 U5427 (.A1(W3229), .A2(I786), .ZN(W5427));
	NANDX1 U5437 (.A1(W3400), .A2(O154), .ZN(W5437));
	NANDX1 U5441 (.A1(W652), .A2(I910), .ZN(O327));
	INVX1 U5467 (.I(W932), .ZN(W5467));
	NANDX1 U5487 (.A1(W3928), .A2(W1036), .ZN(W5487));
	NANDX1 U5502 (.A1(W4305), .A2(W1562), .ZN(O118));
	INVX1 U5503 (.I(W1253), .ZN(O184));
	NOR2X1 U5513 (.A1(W2837), .A2(I4435), .ZN(W5513));
	NANDX1 U5515 (.A1(W4414), .A2(W2718), .ZN(W5515));
	INVX1 U5527 (.I(W3646), .ZN(O260));
	INVX1 U5533 (.I(W4619), .ZN(W5533));
	INVX1 U5546 (.I(W3657), .ZN(W5546));
	INVX1 U5559 (.I(W5197), .ZN(W5559));
	INVX1 U5567 (.I(W5404), .ZN(O225));
	INVX1 U5587 (.I(I1913), .ZN(W5587));
	INVX1 U5602 (.I(I664), .ZN(O389));
	NOR2X1 U5613 (.A1(W3873), .A2(W2725), .ZN(O367));
	NANDX1 U5618 (.A1(W3084), .A2(W935), .ZN(W5618));
	NANDX1 U5638 (.A1(O21), .A2(W4163), .ZN(O5));
	INVX1 U5645 (.I(W3950), .ZN(O452));
	NOR2X1 U5654 (.A1(W2620), .A2(W585), .ZN(O421));
	NANDX1 U5656 (.A1(O365), .A2(I3795), .ZN(O87));
	NANDX1 U5664 (.A1(W2080), .A2(W1913), .ZN(W5664));
	INVX1 U5683 (.I(W2411), .ZN(W5683));
	NOR2X1 U5685 (.A1(W1980), .A2(W2937), .ZN(O310));
	NOR2X1 U5698 (.A1(I2939), .A2(W1659), .ZN(O429));
	NANDX1 U5700 (.A1(W4357), .A2(W470), .ZN(O64));
	NOR2X1 U5709 (.A1(W3629), .A2(W4499), .ZN(W5709));
	NANDX1 U5715 (.A1(W370), .A2(I3406), .ZN(W5715));
	NANDX1 U5730 (.A1(W1425), .A2(W2487), .ZN(W5730));
	NOR2X1 U5743 (.A1(W582), .A2(W284), .ZN(W5743));
	NANDX1 U5753 (.A1(W4139), .A2(I1216), .ZN(O235));
	NANDX1 U5790 (.A1(W3520), .A2(W3799), .ZN(W5790));
	INVX1 U5796 (.I(W5709), .ZN(O170));
	INVX1 U5799 (.I(W5375), .ZN(W5799));
	NANDX1 U5827 (.A1(I1433), .A2(W1339), .ZN(W5827));
	NANDX1 U5846 (.A1(W1774), .A2(W2753), .ZN(W5846));
	NOR2X1 U5866 (.A1(W2789), .A2(W4063), .ZN(O347));
	INVX1 U5873 (.I(I1375), .ZN(O208));
	INVX1 U5886 (.I(W1726), .ZN(W5886));
	NOR2X1 U5894 (.A1(W5467), .A2(W4421), .ZN(O481));
	INVX1 U5911 (.I(W3104), .ZN(W5911));
	NOR2X1 U5922 (.A1(W1153), .A2(W2413), .ZN(W5922));
	NANDX1 U5951 (.A1(W4824), .A2(W3991), .ZN(W5951));
	NOR2X1 U5953 (.A1(W4267), .A2(I3986), .ZN(W5953));
	NOR2X1 U5959 (.A1(O76), .A2(W5356), .ZN(W5959));
	NOR2X1 U5970 (.A1(W3495), .A2(W2984), .ZN(O71));
	INVX1 U5976 (.I(W1416), .ZN(O247));
	INVX1 U5978 (.I(I4872), .ZN(W5978));
	NOR2X1 U5982 (.A1(W4334), .A2(W5336), .ZN(W5982));
	INVX1 U5989 (.I(I4605), .ZN(W5989));
	NANDX1 U5991 (.A1(I4645), .A2(W5117), .ZN(O489));
	INVX1 U5996 (.I(I3014), .ZN(W5996));
	NANDX1 U5999 (.A1(W1251), .A2(W3405), .ZN(W5999));
	NOR2X1 U6010 (.A1(O430), .A2(W3953), .ZN(O412));
	NANDX1 U6018 (.A1(W4831), .A2(O289), .ZN(O308));
	NOR2X1 U6028 (.A1(W1781), .A2(I4117), .ZN(O409));
	NOR2X1 U6035 (.A1(O98), .A2(W3126), .ZN(W6035));
	NOR2X1 U6053 (.A1(I432), .A2(W4607), .ZN(W6053));
	INVX1 U6071 (.I(W5388), .ZN(O90));
	INVX1 U6083 (.I(W1655), .ZN(W6083));
	INVX1 U6086 (.I(W2225), .ZN(W6086));
	NOR2X1 U6087 (.A1(W2745), .A2(W3164), .ZN(W6087));
	INVX1 U6100 (.I(W1353), .ZN(W6100));
	INVX1 U6113 (.I(I1971), .ZN(O461));
	NOR2X1 U6118 (.A1(W2786), .A2(W5054), .ZN(W6118));
	NANDX1 U6145 (.A1(W3663), .A2(W1417), .ZN(W6145));
	NOR2X1 U6173 (.A1(I2802), .A2(W5099), .ZN(W6173));
	NANDX1 U6178 (.A1(W885), .A2(W5978), .ZN(O213));
	NANDX1 U6204 (.A1(O241), .A2(W2349), .ZN(W6204));
	NOR2X1 U6207 (.A1(I1492), .A2(W5799), .ZN(O16));
	INVX1 U6208 (.I(W5333), .ZN(O302));
	INVX1 U6225 (.I(W1519), .ZN(O307));
	INVX1 U6248 (.I(W2040), .ZN(O268));
	INVX1 U6262 (.I(W2974), .ZN(W6262));
	INVX1 U6278 (.I(O71), .ZN(W6278));
	NANDX1 U6291 (.A1(W3852), .A2(W4754), .ZN(O446));
	INVX1 U6292 (.I(I818), .ZN(W6292));
	NOR2X1 U6298 (.A1(W1637), .A2(W6145), .ZN(O313));
	INVX1 U6314 (.I(W674), .ZN(W6314));
	NANDX1 U6320 (.A1(W697), .A2(W3435), .ZN(W6320));
	NANDX1 U6322 (.A1(W3216), .A2(W1672), .ZN(O320));
	INVX1 U6340 (.I(I490), .ZN(O160));
	NOR2X1 U6352 (.A1(W3843), .A2(W3833), .ZN(O232));
	INVX1 U6375 (.I(W568), .ZN(W6375));
	NOR2X1 U6382 (.A1(W5911), .A2(W1211), .ZN(W6382));
	NANDX1 U6383 (.A1(W6100), .A2(W6118), .ZN(W6383));
	NANDX1 U6385 (.A1(W5827), .A2(W304), .ZN(O83));
	NOR2X1 U6386 (.A1(W3227), .A2(W595), .ZN(W6386));
	NOR2X1 U6391 (.A1(W3344), .A2(W1160), .ZN(W6391));
	NOR2X1 U6399 (.A1(W5533), .A2(W5959), .ZN(O24));
	NANDX1 U6402 (.A1(W5378), .A2(W5989), .ZN(O340));
	NOR2X1 U6403 (.A1(W6262), .A2(W2012), .ZN(W6403));
	INVX1 U6406 (.I(I2338), .ZN(W6406));
	INVX1 U6408 (.I(W3036), .ZN(W6408));
	NANDX1 U6411 (.A1(W3430), .A2(W5113), .ZN(O273));
	NOR2X1 U6417 (.A1(W748), .A2(O24), .ZN(W6417));
	INVX1 U6431 (.I(W2247), .ZN(W6431));
	NOR2X1 U6446 (.A1(W5683), .A2(W3699), .ZN(O410));
	INVX1 U6455 (.I(W3991), .ZN(W6455));
	INVX1 U6464 (.I(I4178), .ZN(O301));
	NOR2X1 U6468 (.A1(W53), .A2(I3552), .ZN(O53));
	NOR2X1 U6474 (.A1(W9), .A2(W2427), .ZN(O398));
	NANDX1 U6476 (.A1(W5241), .A2(W4738), .ZN(W6476));
	NOR2X1 U6512 (.A1(W898), .A2(W625), .ZN(W6512));
	NANDX1 U6524 (.A1(I4817), .A2(W4304), .ZN(W6524));
	INVX1 U6529 (.I(W2146), .ZN(O207));
	INVX1 U6533 (.I(W2771), .ZN(W6533));
	NOR2X1 U6559 (.A1(W5922), .A2(W2754), .ZN(W6559));
	NANDX1 U6563 (.A1(I32), .A2(W5153), .ZN(O201));
	INVX1 U6569 (.I(W3301), .ZN(O140));
	NOR2X1 U6572 (.A1(W5013), .A2(I4231), .ZN(W6572));
	NOR2X1 U6579 (.A1(W5587), .A2(I2095), .ZN(O122));
	NOR2X1 U6586 (.A1(W4993), .A2(W3032), .ZN(W6586));
	INVX1 U6594 (.I(W5715), .ZN(W6594));
	NANDX1 U6603 (.A1(W4468), .A2(W6087), .ZN(O451));
	INVX1 U6625 (.I(W204), .ZN(O124));
	NANDX1 U6629 (.A1(W5373), .A2(W1186), .ZN(O40));
	INVX1 U6636 (.I(W4754), .ZN(W6636));
	NOR2X1 U6654 (.A1(W3897), .A2(W4118), .ZN(O233));
	NOR2X1 U6687 (.A1(W5356), .A2(W4435), .ZN(O326));
	INVX1 U6713 (.I(W4517), .ZN(O137));
	NANDX1 U6725 (.A1(W6391), .A2(I2243), .ZN(O392));
	NOR2X1 U6740 (.A1(W5487), .A2(O160), .ZN(W6740));
	INVX1 U6746 (.I(W5036), .ZN(W6746));
	INVX1 U6751 (.I(W4920), .ZN(O175));
	NANDX1 U6765 (.A1(W3878), .A2(I3168), .ZN(W6765));
	NOR2X1 U6782 (.A1(W132), .A2(W4938), .ZN(W6782));
	NOR2X1 U6785 (.A1(I1670), .A2(W1528), .ZN(O48));
	NOR2X1 U6796 (.A1(I3553), .A2(W6455), .ZN(O386));
	NANDX1 U6801 (.A1(W6524), .A2(I1769), .ZN(W6801));
	INVX1 U6807 (.I(W1172), .ZN(W6807));
	NOR2X1 U6820 (.A1(W1620), .A2(I3319), .ZN(W6820));
	NANDX1 U6824 (.A1(W2456), .A2(W6292), .ZN(W6824));
	NOR2X1 U6848 (.A1(W1538), .A2(W2928), .ZN(O345));
	INVX1 U6860 (.I(W3968), .ZN(O370));
	INVX1 U6875 (.I(W4598), .ZN(W6875));
	NANDX1 U6876 (.A1(W4229), .A2(W4572), .ZN(O455));
	NOR2X1 U6877 (.A1(W1963), .A2(W2208), .ZN(O112));
	INVX1 U6889 (.I(W3185), .ZN(O435));
	NOR2X1 U6902 (.A1(W3376), .A2(W649), .ZN(W6902));
	NANDX1 U6921 (.A1(W4991), .A2(I4477), .ZN(O188));
	NANDX1 U6922 (.A1(W6476), .A2(I3094), .ZN(O186));
	NOR2X1 U6944 (.A1(I4286), .A2(W4423), .ZN(O445));
	INVX1 U6953 (.I(I1678), .ZN(W6953));
	NOR2X1 U6957 (.A1(W6403), .A2(W4573), .ZN(W6957));
	INVX1 U6963 (.I(W5999), .ZN(O174));
	NANDX1 U6975 (.A1(W4919), .A2(W4822), .ZN(O135));
	NANDX1 U6987 (.A1(W3734), .A2(W4959), .ZN(W6987));
	INVX1 U6988 (.I(W5559), .ZN(W6988));
	NOR2X1 U6997 (.A1(W5546), .A2(W2683), .ZN(O193));
	NANDX1 U7000 (.A1(W4065), .A2(W6636), .ZN(O405));
	NOR2X1 U7011 (.A1(W1285), .A2(W6824), .ZN(O485));
	NOR2X1 U7012 (.A1(W5437), .A2(W4440), .ZN(O240));
	INVX1 U7023 (.I(W3021), .ZN(W7023));
	NOR2X1 U7025 (.A1(I2718), .A2(W4799), .ZN(O397));
	INVX1 U7042 (.I(W3457), .ZN(W7042));
	NOR2X1 U7105 (.A1(I2248), .A2(W4508), .ZN(O23));
	NOR2X1 U7110 (.A1(W1126), .A2(I4595), .ZN(O33));
	NANDX1 U7127 (.A1(W5211), .A2(O244), .ZN(W7127));
	NANDX1 U7145 (.A1(W3859), .A2(W686), .ZN(W7145));
	NANDX1 U7148 (.A1(W5235), .A2(W6035), .ZN(O164));
	NANDX1 U7152 (.A1(W3317), .A2(W2331), .ZN(O223));
	NOR2X1 U7154 (.A1(I3610), .A2(W6053), .ZN(W7154));
	INVX1 U7180 (.I(W2267), .ZN(O245));
	NANDX1 U7200 (.A1(I3136), .A2(W1482), .ZN(O195));
	NANDX1 U7215 (.A1(W2792), .A2(I223), .ZN(O470));
	NANDX1 U7241 (.A1(O233), .A2(W6953), .ZN(W7241));
	INVX1 U7245 (.I(I4506), .ZN(O440));
	NANDX1 U7248 (.A1(W5334), .A2(W902), .ZN(O103));
	NOR2X1 U7281 (.A1(W5618), .A2(W6382), .ZN(O287));
	INVX1 U7304 (.I(W2786), .ZN(O473));
	NOR2X1 U7347 (.A1(W2697), .A2(I807), .ZN(W7347));
	INVX1 U7351 (.I(W2), .ZN(W7351));
	INVX1 U7353 (.I(W3083), .ZN(O393));
	INVX1 U7357 (.I(W2293), .ZN(O96));
	INVX1 U7358 (.I(W5951), .ZN(O443));
	NOR2X1 U7366 (.A1(W2589), .A2(W4033), .ZN(O56));
	NOR2X1 U7377 (.A1(I2679), .A2(I1971), .ZN(W7377));
	NANDX1 U7381 (.A1(W513), .A2(W7042), .ZN(W7381));
	NANDX1 U7383 (.A1(O411), .A2(W6204), .ZN(O254));
	INVX1 U7407 (.I(W6746), .ZN(O396));
	INVX1 U7433 (.I(I121), .ZN(W7433));
	NOR2X1 U7446 (.A1(W3562), .A2(W4965), .ZN(W7446));
	NOR2X1 U7452 (.A1(W3288), .A2(I187), .ZN(O1));
	NANDX1 U7458 (.A1(W5982), .A2(W6431), .ZN(O494));
	INVX1 U7462 (.I(W441), .ZN(O269));
	INVX1 U7463 (.I(W6572), .ZN(W7463));
	INVX1 U7465 (.I(O318), .ZN(O249));
	NANDX1 U7467 (.A1(W6408), .A2(I3383), .ZN(O41));
	NOR2X1 U7468 (.A1(W4451), .A2(W7145), .ZN(O344));
	NOR2X1 U7499 (.A1(I4495), .A2(W6417), .ZN(O328));
	INVX1 U7517 (.I(W2408), .ZN(O321));
	INVX1 U7519 (.I(I174), .ZN(W7519));
	NANDX1 U7520 (.A1(W5790), .A2(W2498), .ZN(O448));
	NOR2X1 U7529 (.A1(W1292), .A2(W1219), .ZN(W7529));
	NOR2X1 U7543 (.A1(W4597), .A2(W5174), .ZN(O495));
	NANDX1 U7564 (.A1(W2216), .A2(I4749), .ZN(O252));
	NOR2X1 U7570 (.A1(I3137), .A2(W6902), .ZN(O468));
	NANDX1 U7585 (.A1(I3557), .A2(W5996), .ZN(O59));
	NANDX1 U7592 (.A1(I2282), .A2(W4121), .ZN(W7592));
	NOR2X1 U7599 (.A1(W2489), .A2(I2919), .ZN(O11));
	NOR2X1 U7614 (.A1(W5233), .A2(W7592), .ZN(O150));
	NOR2X1 U7678 (.A1(I4847), .A2(W5886), .ZN(W7678));
	NOR2X1 U7680 (.A1(W188), .A2(W1548), .ZN(O361));
	NANDX1 U7700 (.A1(I3330), .A2(W5009), .ZN(O222));
	NANDX1 U7730 (.A1(W428), .A2(W6765), .ZN(O349));
	NOR2X1 U7744 (.A1(W2019), .A2(W4886), .ZN(O50));
	INVX1 U7752 (.I(I4775), .ZN(W7752));
	NANDX1 U7757 (.A1(W2476), .A2(I727), .ZN(O329));
	NANDX1 U7771 (.A1(W4552), .A2(W2604), .ZN(O12));
	NANDX1 U7778 (.A1(W7154), .A2(W3939), .ZN(O382));
	NOR2X1 U7784 (.A1(I3474), .A2(W3591), .ZN(O387));
	NOR2X1 U7787 (.A1(I1249), .A2(W4476), .ZN(O447));
	NANDX1 U7816 (.A1(W5515), .A2(W3288), .ZN(O100));
	NOR2X1 U7833 (.A1(W1564), .A2(W5073), .ZN(O423));
	NANDX1 U7842 (.A1(W1767), .A2(W185), .ZN(O45));
	NOR2X1 U7880 (.A1(W5125), .A2(W3289), .ZN(W7880));
	NANDX1 U7897 (.A1(W2346), .A2(W3215), .ZN(O125));
	NANDX1 U7912 (.A1(O231), .A2(W2327), .ZN(O203));
	INVX1 U7917 (.I(I3001), .ZN(W7917));
	NOR2X1 U7921 (.A1(O447), .A2(W5283), .ZN(O366));
	NOR2X1 U7932 (.A1(W702), .A2(W3037), .ZN(O237));
	NOR2X1 U7946 (.A1(I3680), .A2(W5846), .ZN(O403));
	NOR2X1 U7959 (.A1(I892), .A2(W760), .ZN(W7959));
	INVX1 U7973 (.I(W1610), .ZN(O484));
	INVX1 U7981 (.I(W4966), .ZN(O101));
	NOR2X1 U7993 (.A1(W6278), .A2(W7959), .ZN(O166));
	NOR2X1 U8008 (.A1(W2237), .A2(W5513), .ZN(W8008));
	NOR2X1 U8018 (.A1(W5403), .A2(W1589), .ZN(O284));
	NOR2X1 U8027 (.A1(W1923), .A2(W2183), .ZN(O85));
	NOR2X1 U8057 (.A1(I4449), .A2(W1642), .ZN(O242));
	INVX1 U8069 (.I(W2987), .ZN(O278));
	INVX1 U8081 (.I(W5382), .ZN(O156));
	INVX1 U8095 (.I(I2180), .ZN(W8095));
	INVX1 U8097 (.I(W3278), .ZN(O304));
	NANDX1 U8107 (.A1(W6083), .A2(W5405), .ZN(O374));
	INVX1 U8167 (.I(W4883), .ZN(W8167));
	NOR2X1 U8177 (.A1(W6782), .A2(W3105), .ZN(O36));
	INVX1 U8231 (.I(W4608), .ZN(W8231));
	NANDX1 U8263 (.A1(W1737), .A2(W6512), .ZN(O465));
	INVX1 U8276 (.I(I3298), .ZN(O342));
	NOR2X1 U8324 (.A1(W1821), .A2(W3380), .ZN(O158));
	NOR2X1 U8329 (.A1(O36), .A2(W7241), .ZN(O218));
	NOR2X1 U8351 (.A1(W3127), .A2(I435), .ZN(W8351));
	INVX1 U8360 (.I(W4296), .ZN(O163));
	NANDX1 U8361 (.A1(W6586), .A2(W7377), .ZN(O107));
	INVX1 U8364 (.I(I343), .ZN(O360));
	INVX1 U8400 (.I(W2689), .ZN(O341));
	NOR2X1 U8401 (.A1(W3723), .A2(W6957), .ZN(O28));
	INVX1 U8476 (.I(W6987), .ZN(W8476));
	INVX1 U8478 (.I(W4657), .ZN(O442));
	NOR2X1 U8479 (.A1(W4673), .A2(W7381), .ZN(O95));
	INVX1 U8480 (.I(W7752), .ZN(O78));
	INVX1 U8485 (.I(W7127), .ZN(W8485));
	NOR2X1 U8506 (.A1(W7433), .A2(W6807), .ZN(W8506));
	NOR2X1 U8526 (.A1(W2630), .A2(W6320), .ZN(O343));
	NOR2X1 U8533 (.A1(W2903), .A2(W3265), .ZN(O270));
	NANDX1 U8558 (.A1(I1873), .A2(W6383), .ZN(O264));
	INVX1 U8561 (.I(W6083), .ZN(O214));
	NANDX1 U8569 (.A1(W3237), .A2(W2818), .ZN(O462));
	NANDX1 U8600 (.A1(W8095), .A2(W1311), .ZN(O444));
	NANDX1 U8613 (.A1(W5088), .A2(W5730), .ZN(O82));
	NOR2X1 U8618 (.A1(W5324), .A2(O459), .ZN(O229));
	INVX1 U8633 (.I(W7917), .ZN(O22));
	NOR2X1 U8635 (.A1(I3916), .A2(W5372), .ZN(W8635));
	NANDX1 U8651 (.A1(W5664), .A2(W4035), .ZN(O142));
	NANDX1 U8686 (.A1(W4488), .A2(W8485), .ZN(O102));
	NANDX1 U8702 (.A1(W2194), .A2(O98), .ZN(O331));
	NOR2X1 U8705 (.A1(W6086), .A2(W7347), .ZN(O439));
	INVX1 U8732 (.I(W7446), .ZN(O31));
	INVX1 U8778 (.I(W6875), .ZN(O438));
	INVX1 U8790 (.I(I1788), .ZN(O8));
	NANDX1 U8795 (.A1(W3955), .A2(W3363), .ZN(W8795));
	NANDX1 U8807 (.A1(W6406), .A2(W6375), .ZN(O305));
	INVX1 U8885 (.I(W2416), .ZN(O106));
	INVX1 U8902 (.I(W796), .ZN(O297));
	NOR2X1 U8923 (.A1(W5101), .A2(W8795), .ZN(O432));
	NANDX1 U8927 (.A1(W2497), .A2(W4985), .ZN(O9));
	INVX1 U8934 (.I(W8008), .ZN(O417));
	NANDX1 U8942 (.A1(W2302), .A2(W3052), .ZN(O60));
	NOR2X1 U9008 (.A1(W6386), .A2(W7880), .ZN(O26));
	NANDX1 U9017 (.A1(W2957), .A2(W3810), .ZN(O413));
	NANDX1 U9021 (.A1(W2131), .A2(I3117), .ZN(O492));
	INVX1 U9042 (.I(W4466), .ZN(O425));
	NANDX1 U9051 (.A1(W4947), .A2(W7351), .ZN(O486));
	INVX1 U9059 (.I(W6988), .ZN(O350));
	NOR2X1 U9079 (.A1(W5953), .A2(W4129), .ZN(O337));
	NOR2X1 U9084 (.A1(I412), .A2(I3429), .ZN(O169));
	NANDX1 U9092 (.A1(W6820), .A2(W1763), .ZN(O228));
	NOR2X1 U9118 (.A1(W3247), .A2(W2745), .ZN(W9118));
	NANDX1 U9134 (.A1(W9118), .A2(I2798), .ZN(W9134));
	INVX1 U9151 (.I(W3363), .ZN(O138));
	INVX1 U9213 (.I(W3565), .ZN(W9213));
	NANDX1 U9224 (.A1(W4865), .A2(I1802), .ZN(O496));
	INVX1 U9229 (.I(W8351), .ZN(O493));
	NOR2X1 U9249 (.A1(W3637), .A2(W2513), .ZN(O167));
	INVX1 U9268 (.I(W5363), .ZN(O357));
	NANDX1 U9274 (.A1(I2897), .A2(W7023), .ZN(O70));
	NANDX1 U9290 (.A1(W2331), .A2(W4164), .ZN(O37));
	NOR2X1 U9323 (.A1(W5743), .A2(O263), .ZN(O322));
	INVX1 U9341 (.I(W8476), .ZN(O230));
	INVX1 U9343 (.I(W2547), .ZN(O388));
	NOR2X1 U9364 (.A1(W6533), .A2(I3419), .ZN(O399));
	NOR2X1 U9384 (.A1(W6173), .A2(W4412), .ZN(O38));
	NOR2X1 U9393 (.A1(W3344), .A2(I4573), .ZN(O126));
	NOR2X1 U9407 (.A1(W8231), .A2(W4909), .ZN(O113));
	NANDX1 U9445 (.A1(I3980), .A2(I1350), .ZN(O266));
	NANDX1 U9541 (.A1(W6559), .A2(W4271), .ZN(O20));
	NOR2X1 U9547 (.A1(W9134), .A2(W1026), .ZN(O69));
	INVX1 U9566 (.I(W8167), .ZN(O17));
	NANDX1 U9617 (.A1(W4706), .A2(W1182), .ZN(O110));
	INVX1 U9621 (.I(W8506), .ZN(O404));
	NANDX1 U9719 (.A1(I2746), .A2(I3686), .ZN(O131));
	NOR2X1 U9725 (.A1(W4794), .A2(W6801), .ZN(O375));
	NANDX1 U9756 (.A1(O320), .A2(W6314), .ZN(O89));
	NOR2X1 U9767 (.A1(W6594), .A2(W5073), .ZN(O499));
	NANDX1 U9777 (.A1(I3590), .A2(W322), .ZN(O6));
	NANDX1 U9826 (.A1(W9213), .A2(W6740), .ZN(O290));
	NANDX1 U9841 (.A1(W1720), .A2(W7463), .ZN(O144));
	NANDX1 U9882 (.A1(I1299), .A2(W1067), .ZN(O63));
	NANDX1 U9884 (.A1(W8635), .A2(W5427), .ZN(O295));
	INVX1 U9888 (.I(W4325), .ZN(O251));
	NANDX1 U9898 (.A1(W7678), .A2(W5426), .ZN(O205));
	NANDX1 U9960 (.A1(W7529), .A2(W3452), .ZN(O18));
	INVX1 U9964 (.I(W378), .ZN(O281));
	INVX1 U9976 (.I(W7519), .ZN(O414));
	
endmodule
